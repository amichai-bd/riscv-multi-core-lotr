@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 10 57 73 00 10 00
@000000A8
13 01 01 FE 23 2E 81 00 13 04 01 02 23 26 04 FE
6F 00 00 01 83 27 C4 FE 93 87 17 00 23 26 F4 FE
03 27 C4 FE B7 47 01 00 93 87 F7 87 E3 D4 E7 FE
13 00 00 00 13 00 00 00 03 24 C1 01 13 01 01 02
67 80 00 00 13 01 01 FC 23 2E 81 02 13 04 01 04
23 26 A4 FC 23 24 B4 FC 23 22 C4 FC 83 27 84 FC
93 87 17 14 93 97 17 00 03 27 44 FC B3 07 F7 00
23 22 F4 FE B7 17 00 00 93 87 07 E1 23 20 F4 FE
03 27 C4 FC 93 07 07 00 93 97 27 00 B3 87 E7 00
93 97 47 00 93 87 17 00 23 2E F4 FC 23 26 04 FE
6F 00 40 03 03 27 44 FE 83 27 C4 FE 33 07 F7 40
83 27 04 FE B3 07 F7 00 13 97 27 00 B7 07 40 03
B3 07 F7 00 23 A0 07 00 83 27 C4 FE 93 87 07 05
23 26 F4 FE 03 27 C4 FE B7 17 00 00 93 87 07 96
E3 D2 E7 FC 23 24 04 FE 6F 00 80 03 03 27 44 FE
83 27 84 FE 33 07 F7 40 83 27 04 FE B3 07 F7 00
13 97 27 00 B7 07 40 03 B3 07 F7 00 13 07 F0 FF
23 A0 E7 00 83 27 84 FE 93 87 07 05 23 24 F4 FE
03 27 84 FE 83 27 C4 FD E3 42 F7 FC 13 00 00 00
13 00 00 00 03 24 C1 03 13 01 01 04 67 80 00 00
13 01 01 FD 23 26 81 02 13 04 01 03 23 2E A4 FC
23 2C B4 FC 83 27 C4 FD 83 C7 07 00 A3 07 F4 FE
83 27 84 FD 03 C7 07 00 83 27 C4 FD 23 80 E7 00
83 27 84 FD 03 47 F4 FE 23 80 E7 00 13 00 00 00
03 24 C1 02 13 01 01 03 67 80 00 00 13 01 01 FD
23 26 11 02 23 24 81 02 13 04 01 03 23 2E A4 FC
23 2C B4 FC 23 26 04 FE 6F 00 00 0E 23 24 04 FE
6F 00 40 0B 83 27 84 FE 03 27 C4 FD B3 07 F7 00
03 C7 07 00 83 27 84 FE 93 87 17 00 83 26 C4 FD
B3 87 F6 00 83 C7 07 00 63 F0 E7 08 83 27 84 FE
03 27 C4 FD B3 06 F7 00 83 27 84 FE 93 87 17 00
03 27 C4 FD B3 07 F7 00 93 85 07 00 13 85 06 00
EF F0 1F F4 83 27 84 FE 03 27 C4 FD B3 07 F7 00
83 C7 07 00 13 06 80 02 83 25 84 FE 13 85 07 00
EF F0 5F E2 83 27 84 FE 93 87 17 00 03 27 C4 FD
B3 07 F7 00 83 C7 07 00 13 87 07 00 83 27 84 FE
93 87 17 00 13 06 80 02 93 85 07 00 13 05 07 00
EF F0 5F DF EF F0 DF DA 83 27 84 FE 93 87 17 00
23 24 F4 FE 03 27 84 FD 83 27 C4 FE B3 07 F7 40
93 87 F7 FF 03 27 84 FE E3 4E F7 F2 83 27 C4 FE
93 87 17 00 23 26 F4 FE 83 27 84 FD 93 87 F7 FF
03 27 C4 FE E3 4C F7 F0 13 00 00 00 13 00 00 00
83 20 C1 02 03 24 81 02 13 01 01 03 67 80 00 00
13 01 01 FD 23 26 11 02 23 24 81 02 13 04 01 03
23 2E A4 FC 93 87 05 00 13 07 06 00 A3 0D F4 FC
93 07 07 00 23 0D F4 FC 83 47 A4 FD 03 27 C4 FD
B3 07 F7 00 83 C7 07 00 A3 03 F4 FE 83 47 B4 FD
93 87 F7 FF A3 07 F4 FE 83 47 B4 FD 23 24 F4 FE
6F 00 80 0C 83 27 84 FE 03 27 C4 FD B3 07 F7 00
83 C7 07 00 03 47 74 FE 63 62 F7 0A 83 47 F4 FE
93 87 17 00 A3 07 F4 FE 83 47 F4 FE 03 27 C4 FD
B3 06 F7 00 83 27 84 FE 03 27 C4 FD B3 07 F7 00
93 85 07 00 13 85 06 00 EF F0 9F DF 83 47 F4 FE
03 27 C4 FD B3 07 F7 00 83 C7 07 00 13 87 07 00
83 47 F4 FE 13 06 00 00 93 85 07 00 13 05 07 00
EF F0 5F CD 83 27 84 FE 03 27 C4 FD B3 07 F7 00
83 C7 07 00 13 06 00 00 83 25 84 FE 13 85 07 00
EF F0 5F CB 83 47 F4 FE 03 27 C4 FD B3 07 F7 00
03 C7 07 00 83 27 84 FE 83 26 C4 FD B3 87 F6 00
83 C7 07 00 63 04 F7 00 EF F0 9F C4 83 27 84 FE
93 87 17 00 23 24 F4 FE 83 47 A4 FD 03 27 84 FE
E3 4A F7 F2 83 47 F4 FE 93 87 17 00 03 27 C4 FD
B3 06 F7 00 83 47 A4 FD 03 27 C4 FD B3 07 F7 00
93 85 07 00 13 85 06 00 EF F0 9F D4 83 47 F4 FE
93 87 17 00 03 27 C4 FD B3 07 F7 00 83 C7 07 00
13 87 07 00 83 47 F4 FE 93 87 17 00 13 06 00 00
93 85 07 00 13 05 07 00 EF F0 DF C1 83 47 A4 FD
03 27 C4 FD B3 07 F7 00 83 C7 07 00 13 87 07 00
83 47 A4 FD 13 06 00 00 93 85 07 00 13 05 07 00
EF F0 5F BF 83 47 F4 FE 93 87 17 00 03 27 C4 FD
B3 07 F7 00 03 C7 07 00 83 47 A4 FD 83 26 C4 FD
B3 87 F6 00 83 C7 07 00 63 04 F7 00 EF F0 5F B8
83 47 F4 FE 93 87 17 00 13 85 07 00 83 20 C1 02
03 24 81 02 13 01 01 03 67 80 00 00 13 01 01 FD
23 26 11 02 23 24 81 02 23 22 91 02 13 04 01 03
23 2E A4 FC 93 86 05 00 A3 0D D4 FC 93 06 06 00
23 0D D4 FC 93 06 01 00 93 84 06 00 03 46 A4 FD
83 46 B4 FD B3 06 D6 40 93 86 16 00 13 86 F6 FF
23 24 C4 FE 13 86 06 00 13 0E 06 00 93 0E 00 00
13 56 DE 01 93 98 3E 00 B3 68 16 01 13 18 3E 00
13 86 06 00 13 03 06 00 93 03 00 00 13 56 D3 01
93 97 33 00 B3 67 F6 00 13 17 33 00 93 87 06 00
93 87 F7 00 93 D7 47 00 93 97 47 00 33 01 F1 40
93 07 01 00 93 87 07 00 23 22 F4 FE 93 07 F0 FF
23 26 F4 FE 83 27 C4 FE 93 87 17 00 23 26 F4 FE
03 27 44 FE 83 27 C4 FE B3 07 F7 00 03 47 B4 FD
23 80 E7 00 83 27 C4 FE 93 87 17 00 23 26 F4 FE
03 27 44 FE 83 27 C4 FE B3 07 F7 00 03 47 A4 FD
23 80 E7 00 6F 00 C0 10 83 27 C4 FE 13 87 F7 FF
23 26 E4 FE 03 27 44 FE B3 07 F7 00 83 C7 07 00
23 0D F4 FC 83 27 C4 FE 13 87 F7 FF 23 26 E4 FE
03 27 44 FE B3 07 F7 00 83 C7 07 00 A3 0D F4 FC
03 47 A4 FD 83 47 B4 FD 13 06 07 00 93 85 07 00
03 25 C4 FD EF F0 DF CD 93 07 05 00 A3 01 F4 FE
83 47 34 FE 13 87 F7 FF 83 47 B4 FD 63 D6 E7 04
83 27 C4 FE 93 87 17 00 23 26 F4 FE 03 27 44 FE
83 27 C4 FE B3 07 F7 00 03 47 B4 FD 23 80 E7 00
83 27 C4 FE 93 87 17 00 23 26 F4 FE 83 47 34 FE
93 87 F7 FF 13 F7 F7 0F 83 26 44 FE 83 27 C4 FE
B3 87 F6 00 23 80 E7 00 83 47 34 FE 13 87 17 00
83 47 A4 FD 63 56 F7 04 83 27 C4 FE 93 87 17 00
23 26 F4 FE 83 47 34 FE 93 87 17 00 13 F7 F7 0F
83 26 44 FE 83 27 C4 FE B3 87 F6 00 23 80 E7 00
83 27 C4 FE 93 87 17 00 23 26 F4 FE 03 27 44 FE
83 27 C4 FE B3 07 F7 00 03 47 A4 FD 23 80 E7 00
83 27 C4 FE E3 DA 07 EE 13 81 04 00 13 00 00 00
13 01 04 FD 83 20 C1 02 03 24 81 02 83 24 41 02
13 01 01 03 67 80 00 00 13 01 01 FE 23 2E 81 00
13 04 01 02 23 26 A4 FE 23 24 B4 FE 03 27 C4 FE
83 27 84 FE 63 54 F7 00 93 07 07 00 13 85 07 00
03 24 C1 01 13 01 01 02 67 80 00 00 13 01 01 FD
23 26 11 02 23 24 81 02 13 04 01 03 23 2E A4 FC
23 2C B4 FC 93 07 10 00 23 26 F4 FE 6F 00 80 0B
23 24 04 FE 6F 00 40 09 03 27 84 FE 83 27 C4 FE
B3 07 F7 00 13 87 F7 FF 83 27 84 FD 93 87 F7 FF
93 85 07 00 13 05 07 00 EF F0 1F F8 23 22 A4 FE
83 27 C4 FE 13 97 17 00 83 27 84 FE B3 07 F7 00
13 87 F7 FF 83 27 84 FD 93 87 F7 FF 93 85 07 00
13 05 07 00 EF F0 5F F5 23 20 A4 FE 83 27 84 FE
93 F7 F7 0F 03 27 44 FE 13 77 F7 0F 83 26 04 FE
93 F6 F6 0F 13 06 07 00 93 85 07 00 03 25 C4 FD
EF 00 80 05 83 27 C4 FE 93 97 17 00 03 27 84 FE
B3 07 F7 00 23 24 F4 FE 83 27 84 FD 93 87 F7 FF
03 27 84 FE E3 42 F7 F6 83 27 C4 FE 93 97 17 00
23 26 F4 FE 03 27 84 FD 83 27 C4 FE E3 C2 E7 F4
13 00 00 00 13 00 00 00 83 20 C1 02 03 24 81 02
13 01 01 03 67 80 00 00 13 01 01 FA 23 2E 11 04
23 2C 81 04 23 2A 91 04 23 28 21 05 23 26 31 05
23 24 41 05 23 22 51 05 23 20 61 05 23 2E 71 03
13 04 01 06 23 26 A4 FA 13 85 05 00 93 05 06 00
13 86 06 00 93 06 05 00 A3 05 D4 FA 93 86 05 00
23 05 D4 FA 93 06 06 00 A3 04 D4 FA 93 06 01 00
93 84 06 00 03 46 A4 FA 83 46 B4 FA B3 06 D6 40
93 F6 F6 0F 93 86 16 00 23 06 D4 FC 03 46 94 FA
83 46 A4 FA B3 06 D6 40 A3 05 D4 FC 83 46 C4 FC
13 86 06 00 13 06 F6 FF 23 22 C4 FC 13 8B 06 00
93 0B 00 00 13 56 DB 01 93 9E 3B 00 B3 6E D6 01
13 1E 3B 00 13 8A 06 00 93 0A 00 00 13 56 DA 01
93 93 3A 00 B3 63 76 00 13 13 3A 00 93 86 F6 00
93 D6 46 00 93 96 46 00 33 01 D1 40 93 06 01 00
93 86 06 00 23 20 D4 FC 83 46 B4 FC 13 86 06 00
13 06 F6 FF 23 2E C4 FA 13 89 06 00 93 09 00 00
13 56 D9 01 93 98 39 00 B3 68 16 01 13 18 39 00
13 8F 06 00 93 0F 00 00 13 56 DF 01 93 97 3F 00
B3 67 F6 00 13 17 3F 00 93 87 06 00 93 87 F7 00
93 D7 47 00 93 97 47 00 33 01 F1 40 93 07 01 00
93 87 07 00 23 2C F4 FA A3 06 04 FC 6F 00 C0 03
03 47 B4 FA 83 47 D4 FC B3 07 F7 00 13 87 07 00
83 27 C4 FA 33 87 E7 00 83 47 D4 FC 03 47 07 00
83 26 04 FC B3 87 F6 00 23 80 E7 00 83 47 D4 FC
93 87 17 00 A3 06 F4 FC 03 47 D4 FC 83 47 C4 FC
E3 60 F7 FC 23 07 04 FC 6F 00 00 04 83 47 A4 FA
13 87 17 00 83 47 E4 FC B3 07 F7 00 13 87 07 00
83 27 C4 FA 33 87 E7 00 83 47 E4 FC 03 47 07 00
83 26 84 FB B3 87 F6 00 23 80 E7 00 83 47 E4 FC
93 87 17 00 23 07 F4 FC 03 47 E4 FC 83 47 B4 FC
E3 6E F7 FA A3 06 04 FC 23 07 04 FC 83 47 B4 FA
A3 07 F4 FC 6F 00 00 0F 83 47 D4 FC 03 27 04 FC
B3 07 F7 00 03 C7 07 00 83 47 E4 FC 83 26 84 FB
B3 87 F6 00 83 C7 07 00 63 E2 E7 06 03 47 D4 FC
83 47 F4 FC 83 26 C4 FA B3 87 F6 00 83 26 04 FC
33 87 E6 00 03 47 07 00 23 80 E7 00 83 47 F4 FC
03 27 C4 FA B3 07 F7 00 83 C7 07 00 93 86 07 00
03 47 F4 FC B7 17 00 00 13 86 07 2C 93 05 07 00
13 85 06 00 EF F0 0F E0 EF F0 8F DB 83 47 D4 FC
93 87 17 00 A3 06 F4 FC 6F 00 00 06 03 47 E4 FC
83 47 F4 FC 83 26 C4 FA B3 87 F6 00 83 26 84 FB
33 87 E6 00 03 47 07 00 23 80 E7 00 83 47 F4 FC
03 27 C4 FA B3 07 F7 00 83 C7 07 00 93 86 07 00
03 47 F4 FC B7 17 00 00 13 86 07 2C 93 05 07 00
13 85 06 00 EF F0 0F DA EF F0 8F D5 83 47 E4 FC
93 87 17 00 23 07 F4 FC 83 47 F4 FC 93 87 17 00
A3 07 F4 FC 03 47 D4 FC 83 47 C4 FC 63 7E F7 06
03 47 E4 FC 83 47 B4 FC E3 60 F7 F0 6F 00 C0 06
03 47 D4 FC 83 47 F4 FC 83 26 C4 FA B3 87 F6 00
83 26 04 FC 33 87 E6 00 03 47 07 00 23 80 E7 00
83 47 F4 FC 03 27 C4 FA B3 07 F7 00 83 C7 07 00
93 86 07 00 03 47 F4 FC B7 17 00 00 13 86 07 2C
93 05 07 00 13 85 06 00 EF F0 CF D1 EF F0 4F CD
83 47 D4 FC 93 87 17 00 A3 06 F4 FC 83 47 F4 FC
93 87 17 00 A3 07 F4 FC 03 47 D4 FC 83 47 C4 FC
E3 68 F7 F8 6F 00 C0 06 03 47 E4 FC 83 47 F4 FC
83 26 C4 FA B3 87 F6 00 83 26 84 FB 33 87 E6 00
03 47 07 00 23 80 E7 00 83 47 F4 FC 03 27 C4 FA
B3 07 F7 00 83 C7 07 00 93 86 07 00 03 47 F4 FC
B7 17 00 00 13 86 07 2C 93 05 07 00 13 85 06 00
EF F0 4F CA EF F0 CF C5 83 47 E4 FC 93 87 17 00
23 07 F4 FC 83 47 F4 FC 93 87 17 00 A3 07 F4 FC
03 47 E4 FC 83 47 B4 FC E3 68 F7 F8 13 81 04 00
13 00 00 00 13 01 04 FA 83 20 C1 05 03 24 81 05
83 24 41 05 03 29 01 05 83 29 C1 04 03 2A 81 04
83 2A 41 04 03 2B 01 04 83 2B C1 03 13 01 01 06
67 80 00 00 13 01 01 FD 23 26 11 02 23 24 81 02
13 04 01 03 23 2E A4 FC 23 2C B4 FC 93 07 10 00
23 26 F4 FE 6F 00 00 12 83 27 C4 FE 93 97 27 00
03 27 C4 FD B3 07 F7 00 83 A7 07 00 23 22 F4 FE
83 27 C4 FE 93 87 F7 FF 23 24 F4 FE 6F 00 40 07
83 27 84 FE 93 97 27 00 03 27 C4 FD 33 07 F7 00
83 27 84 FE 93 87 17 00 93 97 27 00 83 26 C4 FD
B3 87 F6 00 03 27 07 00 23 A0 E7 00 83 27 84 FE
93 87 17 00 93 97 27 00 03 27 C4 FD B3 07 F7 00
03 A7 07 00 83 27 84 FE 93 86 17 00 B7 17 00 00
13 86 87 2E 93 85 06 00 13 05 07 00 EF F0 8F B9
EF F0 0F B5 83 27 84 FE 93 87 F7 FF 23 24 F4 FE
83 27 84 FE 63 C0 07 02 83 27 84 FE 93 97 27 00
03 27 C4 FD B3 07 F7 00 83 A7 07 00 03 27 44 FE
E3 48 F7 F6 83 27 84 FE 93 87 17 00 93 97 27 00
03 27 C4 FD B3 07 F7 00 03 27 44 FE 23 A0 E7 00
83 27 84 FE 93 87 17 00 93 97 27 00 03 27 C4 FD
B3 07 F7 00 03 A7 07 00 83 27 84 FE 93 86 17 00
B7 17 00 00 13 86 87 2E 93 85 06 00 13 05 07 00
EF F0 4F B1 EF F0 CF AC 83 27 C4 FE 93 87 17 00
23 26 F4 FE 03 27 C4 FE 83 27 84 FD E3 4E F7 EC
13 00 00 00 13 00 00 00 83 20 C1 02 03 24 81 02
13 01 01 03 67 80 00 00 13 01 01 F4 23 2E 11 0A
23 2C 81 0A 13 04 01 0C B7 07 C0 00 83 A7 07 00
23 2C F4 FC 03 27 84 FD 93 07 70 00 63 0C F7 32
03 27 84 FD 93 07 70 00 63 C6 E7 3C 03 27 84 FD
93 07 60 00 63 06 F7 16 03 27 84 FD 93 07 60 00
63 CA E7 3A 03 27 84 FD 93 07 40 00 63 0A F7 00
03 27 84 FD 93 07 50 00 63 0A F7 0A 6F 00 80 39
EF F0 0F A3 B7 07 40 00 93 87 07 00 83 A5 07 00
03 A6 47 00 83 A6 87 00 03 A7 C7 00 23 2A B4 FA
23 2C C4 FA 23 2E D4 FA 23 20 E4 FC 83 D7 07 01
23 12 F4 FC 93 07 20 01 23 24 F4 FC 23 24 04 FE
6F 00 00 03 83 27 84 FE 13 07 04 FF B3 07 F7 00
83 C7 47 FC 13 06 00 00 83 25 84 FE 13 85 07 00
EF F0 4F A1 83 27 84 FE 93 87 17 00 23 24 F4 FE
03 27 84 FE 83 27 84 FC E3 46 F7 FC EF F0 4F 9B
83 27 84 FC 93 F7 F7 0F 93 87 F7 FF 13 F7 F7 0F
93 07 44 FB 13 06 07 00 93 05 00 00 13 85 07 00
EF F0 CF E2 EF F0 CF 98 6F F0 9F F5 EF F0 4F 98
B7 07 40 00 13 87 47 01 93 07 44 F4 93 06 07 00
13 07 80 04 13 06 07 00 93 85 06 00 13 85 07 00
EF 00 80 2C 93 07 20 01 23 26 F4 FC 23 22 04 FE
6F 00 80 03 83 27 44 FE 93 97 27 00 13 07 04 FF
B3 07 F7 00 03 A7 47 F5 B7 17 00 00 13 86 87 2E
83 25 44 FE 13 05 07 00 EF F0 CF 96 83 27 44 FE
93 87 17 00 23 22 F4 FE 03 27 44 FE 83 27 C4 FC
E3 42 F7 FC EF F0 CF 90 93 07 44 F4 83 25 C4 FC
13 85 07 00 EF F0 1F D0 EF F0 8F 8F 6F F0 1F F7
23 26 04 FE 6F 00 C0 06 83 27 C4 FE 13 97 27 00
B7 07 40 03 B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
03 27 C4 FE B7 17 00 00 93 87 07 2C B3 07 F7 00
13 97 27 00 B7 07 40 03 93 87 07 EC B3 07 F7 00
13 07 F0 FF 23 A0 E7 00 83 27 C4 FE 13 97 27 00
B7 97 40 03 93 87 07 4C B3 07 F7 00 13 07 F0 FF
23 A0 E7 00 83 27 C4 FE 93 87 17 00 23 26 F4 FE
03 27 C4 FE 93 07 F0 04 E3 D8 E7 F8 23 26 04 FE
6F 00 00 09 03 27 C4 FE 93 07 07 00 93 97 27 00
B3 87 E7 00 93 97 67 00 13 87 07 00 B7 07 40 03
B3 07 F7 00 13 07 F0 FF 23 A0 E7 00 03 27 C4 FE
93 07 07 00 93 97 27 00 B3 87 E7 00 93 97 67 00
13 87 07 00 B7 07 40 03 93 87 C7 09 B3 07 F7 00
13 07 F0 FF 23 A0 E7 00 03 27 C4 FE 93 07 07 00
93 97 27 00 B3 87 E7 00 93 97 67 00 13 87 07 00
B7 07 40 03 93 87 C7 13 B3 07 F7 00 13 07 F0 FF
23 A0 E7 00 83 27 C4 FE 93 87 17 00 23 26 F4 FE
03 27 C4 FE 93 07 70 07 E3 D6 E7 F6 EF E0 5F FD
B7 07 40 00 93 87 07 00 83 A5 07 00 03 A6 47 00
83 A6 87 00 03 A7 C7 00 23 20 B4 FA 23 22 C4 FA
23 24 D4 FA 23 26 E4 FA 83 D7 07 01 23 18 F4 FA
93 07 20 01 23 28 F4 FC 23 20 04 FE 6F 00 00 03
83 27 04 FE 13 07 04 FF B3 07 F7 00 83 C7 07 FB
13 06 80 02 83 25 04 FE 13 85 07 00 EF E0 9F FB
83 27 04 FE 93 87 17 00 23 20 F4 FE 03 27 04 FE
83 27 04 FD E3 46 F7 FC EF E0 9F F5 93 07 04 FA
83 25 04 FD 13 85 07 00 EF F0 4F 8D EF E0 5F F4
6F F0 DF F6 EF E0 DF F3 B7 07 40 00 93 87 07 00
83 A5 07 00 03 A6 47 00 83 A6 87 00 03 A7 C7 00
23 26 B4 F8 23 28 C4 F8 23 2A D4 F8 23 2C E4 F8
83 D7 07 01 23 1E F4 F8 93 07 20 01 23 2A F4 FC
23 2E 04 FC 6F 00 80 03 83 27 C4 FD 13 07 04 FF
B3 07 F7 00 83 C7 C7 F9 13 87 07 00 B7 17 00 00
13 86 07 2C 83 25 C4 FD 13 05 07 00 EF E0 9F F1
83 27 C4 FD 93 87 17 00 23 2E F4 FC 03 27 C4 FD
83 27 44 FD E3 42 F7 FC EF E0 9F EB 93 07 C4 F8
83 25 44 FD 13 85 07 00 EF F0 4F D9 EF E0 5F EA
6F F0 5F F6 6F 00 00 00 B3 C7 A5 00 93 F7 37 00
B3 08 C5 00 63 96 07 06 93 07 30 00 63 F2 C7 06
93 77 35 00 13 07 05 00 63 9A 07 0C 13 F6 C8 FF
B3 06 E6 40 93 07 00 02 93 02 00 02 63 C2 D7 06
93 86 05 00 93 07 07 00 63 78 C7 02 03 A8 06 00
93 87 47 00 93 86 46 00 23 AE 07 FF E3 E8 C7 FE
93 07 F6 FF B3 87 E7 40 93 F7 C7 FF 93 87 47 00
33 07 F7 00 B3 85 F5 00 63 68 17 01 67 80 00 00
13 07 05 00 E3 7C 15 FF 83 C7 05 00 13 07 17 00
93 85 15 00 A3 0F F7 FE E3 68 17 FF 67 80 00 00
83 A6 45 00 83 A7 C5 01 83 AF 05 00 03 AF 85 00
83 AE C5 00 03 AE 05 01 03 A3 45 01 03 A8 85 01
23 22 D7 00 83 A6 05 02 23 20 F7 01 23 24 E7 01
23 26 D7 01 23 28 C7 01 23 2A 67 00 23 2C 07 01
23 2E F7 00 13 07 47 02 B3 07 E6 40 23 2E D7 FE
93 85 45 02 E3 C6 F2 FA 6F F0 9F F4 83 C6 05 00
13 07 17 00 93 77 37 00 A3 0F D7 FE 93 85 15 00
E3 8E 07 F0 83 C6 05 00 13 07 17 00 93 77 37 00
A3 0F D7 FE 93 85 15 00 E3 9A 07 FC 6F F0 1F F0
