define DE10_LITE