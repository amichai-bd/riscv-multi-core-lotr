@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
93 00 00 00 13 01 00 00 93 01 00 00 13 02 00 00
93 02 00 00 13 03 00 00 93 03 00 00 13 04 00 00
93 04 00 00 13 05 00 00 93 05 00 00 13 06 00 00
93 06 00 00 13 07 00 00 93 07 00 00 13 88 00 00
93 08 00 00 13 09 00 00 93 09 00 00 13 0A 00 00
93 0A 00 00 13 0B 00 00 93 0B 00 00 13 0C 00 00
93 0C 00 00 13 0D 00 00 93 0D 00 00 13 0E 00 00
93 0E 00 00 13 0F 00 00 93 0F 00 00 B7 00 40 00
37 01 03 04 13 01 11 20 B7 D1 E0 F0 93 81 01 0B
37 02 40 00 13 02 42 00 23 A0 20 00 03 A5 00 00
83 95 00 00 03 86 00 00 83 D6 00 00 03 C7 00 00
23 20 A2 00 23 22 B2 00 23 24 C2 00 23 26 D2 00
23 28 E2 00 83 95 10 00 03 86 10 00 83 D6 10 00
03 C7 10 00 23 2A B2 00 23 2C C2 00 23 2E D2 00
23 20 E2 02 83 95 20 00 03 86 20 00 83 D6 20 00
03 C7 20 00 23 22 B2 02 23 24 C2 02 23 26 D2 02
23 28 E2 02 83 95 30 00 03 86 30 00 83 D6 30 00
03 C7 30 00 23 2A B2 02 23 2C C2 02 23 2E D2 02
23 20 E2 04 B7 C0 AD DE 93 80 F0 EE 37 01 40 00
13 01 81 04 23 00 11 00 A3 00 11 00 23 01 11 00
A3 01 11 00 B7 01 40 00 93 81 C1 04 23 90 11 00
23 91 11 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 73 00 10 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00
