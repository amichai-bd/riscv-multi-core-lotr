@00400800
00 00 C0 3F CD CC 0C 40 BC 08 00 00 48 09 00 00
C8 08 00 00 48 09 00 00 38 09 00 00 48 09 00 00
C8 08 00 00 BC 08 00 00 BC 08 00 00 38 09 00 00
C8 08 00 00 98 08 00 00 98 08 00 00 98 08 00 00
D0 08 00 00 A8 0B 00 00 A8 0B 00 00 CC 0B 00 00
A0 0B 00 00 A0 0B 00 00 34 0C 00 00 CC 0B 00 00
A0 0B 00 00 34 0C 00 00 A0 0B 00 00 CC 0B 00 00
9C 0B 00 00 9C 0B 00 00 9C 0B 00 00 34 0C 00 00
00 01 02 02 03 03 03 03 04 04 04 04 04 04 04 04
05 05 05 05 05 05 05 05 05 05 05 05 05 05 05 05
06 06 06 06 06 06 06 06 06 06 06 06 06 06 06 06
06 06 06 06 06 06 06 06 06 06 06 06 06 06 06 06
07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07
07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07
07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07
07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
