@00400800
