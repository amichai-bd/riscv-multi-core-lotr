@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 C0 1A 73 00 10 00
@000000A8
13 01 01 FD 23 26 11 02 23 24 81 02 23 22 91 02
13 04 01 03 23 2E A4 FC 23 2C B4 FC 23 2A C4 FC
23 26 04 FE 6F 00 80 15 23 24 04 FE 6F 00 80 13
03 27 C4 FE 93 07 07 00 93 97 17 00 B3 87 E7 00
93 97 27 00 13 87 07 00 83 27 44 FD 33 87 E7 00
83 27 84 FE 93 97 27 00 B3 07 F7 00 23 A0 07 00
23 22 04 FE 6F 00 80 0E 03 27 C4 FE 93 07 07 00
93 97 17 00 B3 87 E7 00 93 97 27 00 13 87 07 00
83 27 44 FD 33 87 E7 00 83 27 84 FE 93 97 27 00
B3 07 F7 00 83 A4 07 00 03 27 C4 FE 93 07 07 00
93 97 17 00 B3 87 E7 00 93 97 27 00 13 87 07 00
83 27 C4 FD 33 87 E7 00 83 27 44 FE 93 97 27 00
B3 07 F7 00 83 A6 07 00 03 27 44 FE 93 07 07 00
93 97 17 00 B3 87 E7 00 93 97 27 00 13 87 07 00
83 27 84 FD 33 87 E7 00 83 27 84 FE 93 97 27 00
B3 07 F7 00 83 A7 07 00 93 85 07 00 13 85 06 00
EF 00 40 20 93 07 05 00 13 86 07 00 03 27 C4 FE
93 07 07 00 93 97 17 00 B3 87 E7 00 93 97 27 00
13 87 07 00 83 27 44 FD B3 86 E7 00 33 87 C4 00
83 27 84 FE 93 97 27 00 B3 87 F6 00 23 A0 E7 00
83 27 44 FE 93 87 17 00 23 22 F4 FE 03 27 44 FE
93 07 20 00 E3 DA E7 F0 83 27 84 FE 93 87 17 00
23 24 F4 FE 03 27 84 FE 93 07 20 00 E3 D2 E7 EC
83 27 C4 FE 93 87 17 00 23 26 F4 FE 03 27 C4 FE
93 07 20 00 E3 D2 E7 EA 13 00 00 00 13 00 00 00
83 20 C1 02 03 24 81 02 83 24 41 02 13 01 01 03
67 80 00 00 13 01 01 F7 23 26 11 08 23 24 81 08
13 04 01 09 23 22 04 FE 93 07 10 00 23 20 F4 FC
93 07 20 00 23 22 F4 FC 93 07 30 00 23 24 F4 FC
93 07 40 00 23 26 F4 FC 93 07 50 00 23 28 F4 FC
93 07 60 00 23 2A F4 FC 93 07 70 00 23 2C F4 FC
93 07 80 00 23 2E F4 FC 93 07 90 00 23 20 F4 FE
93 07 90 00 23 2E F4 F8 93 07 80 00 23 20 F4 FA
93 07 70 00 23 22 F4 FA 93 07 60 00 23 24 F4 FA
93 07 50 00 23 26 F4 FA 93 07 40 00 23 28 F4 FA
93 07 30 00 23 2A F4 FA 93 07 20 00 23 2C F4 FA
93 07 10 00 23 2E F4 FA 93 06 84 F7 13 07 C4 F9
93 07 04 FC 13 86 06 00 93 05 07 00 13 85 07 00
EF F0 1F DA 23 26 04 FE 6F 00 80 07 23 24 04 FE
6F 00 80 05 83 27 44 FE 13 87 17 00 23 22 E4 FE
13 97 27 00 B7 17 40 00 93 87 07 F0 B3 06 F7 00
03 27 C4 FE 93 07 07 00 93 97 17 00 B3 87 E7 00
03 27 84 FE B3 87 E7 00 93 97 27 00 93 87 07 FF
B3 87 87 00 83 A7 87 F8 23 A0 F6 00 83 27 84 FE
93 87 17 00 23 24 F4 FE 03 27 84 FE 93 07 20 00
E3 D2 E7 FA 83 27 C4 FE 93 87 17 00 23 26 F4 FE
03 27 C4 FE 93 07 20 00 E3 D2 E7 F8 93 07 00 00
13 85 07 00 83 20 C1 08 03 24 81 08 13 01 01 09
67 80 00 00 13 06 05 00 13 05 00 00 93 F6 15 00
63 84 06 00 33 05 C5 00 93 D5 15 00 13 16 16 00
E3 96 05 FE 67 80 00 00
