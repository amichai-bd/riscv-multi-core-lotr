/*
 User transfer handler FSM 
 Wishbone master unit to 
 handle user transfers 
 between uart host(PC) and device lotr
 */

`timescale 1ns/1ns

module transfer_handler_engine
  #()
   (
    input logic clk,
    input logic rstn,
    input logic interrupt,
    wishbone.master wb_master
    );

endmodule // handshake

   
