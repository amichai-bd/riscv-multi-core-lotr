@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 40 58 73 00 10 00
@000000A8
13 01 01 FD 23 26 81 02 13 04 01 03 93 07 05 00
23 2C B4 FC 23 2A C4 FC A3 0F F4 FC 03 27 84 FD
93 07 07 00 93 97 27 00 B3 87 E7 00 93 97 67 00
23 26 F4 FE 83 27 44 FD 93 97 27 00 23 24 F4 FE
03 27 84 FE 83 27 C4 FE 33 07 F7 00 B7 07 40 03
B3 07 F7 00 23 22 F4 FE 03 27 84 FE 83 27 C4 FE
33 07 F7 00 B7 07 40 03 93 87 07 14 B3 07 F7 00
23 20 F4 FE 83 47 F4 FD 37 07 40 00 13 07 47 09
93 97 27 00 B3 07 F7 00 83 A7 07 00 13 87 07 00
83 27 44 FE 23 A0 E7 00 83 47 F4 FD 37 07 40 00
13 07 87 21 93 97 27 00 B3 07 F7 00 83 A7 07 00
13 87 07 00 83 27 04 FE 23 A0 E7 00 13 00 00 00
03 24 C1 02 13 01 01 03 67 80 00 00 13 01 01 FD
23 26 11 02 23 24 81 02 13 04 01 03 23 2E A4 FC
23 26 04 FE 23 24 04 FE 23 22 04 FE B7 07 C0 00
93 87 07 22 83 A7 07 00 23 22 F4 FE B7 07 C0 00
93 87 47 23 83 A7 07 00 23 24 F4 FE 6F 00 80 0B
83 27 C4 FE 03 27 C4 FD B3 07 F7 00 03 C7 07 00
93 07 A0 00 63 1A F7 02 23 22 04 FE 83 27 84 FE
93 87 27 00 23 24 F4 FE 03 27 84 FE 93 07 80 07
63 14 F7 00 23 24 04 FE 83 27 C4 FE 93 87 17 00
23 26 F4 FE 6F 00 00 07 83 27 C4 FE 03 27 C4 FD
B3 07 F7 00 83 C7 07 00 03 27 84 FE 83 26 44 FE
13 86 06 00 93 05 07 00 13 85 07 00 EF F0 5F E8
83 27 44 FE 93 87 17 00 23 22 F4 FE 03 27 44 FE
93 07 00 05 63 12 F7 02 23 22 04 FE 83 27 84 FE
93 87 27 00 23 24 F4 FE 03 27 84 FE 93 07 80 07
63 14 F7 00 23 24 04 FE 83 27 C4 FE 93 87 17 00
23 26 F4 FE 83 27 C4 FE 03 27 C4 FD B3 07 F7 00
83 C7 07 00 E3 9E 07 F2 B7 07 C0 00 93 87 07 22
03 27 44 FE 23 A0 E7 00 B7 07 C0 00 93 87 47 23
03 27 84 FE 23 A0 E7 00 13 00 00 00 83 20 C1 02
03 24 81 02 13 01 01 03 67 80 00 00 13 01 01 FD
23 26 81 02 13 04 01 03 23 2E A4 FC 23 2C B4 FC
23 2A C4 FC 03 27 84 FD 93 07 07 00 93 97 27 00
B3 87 E7 00 93 97 67 00 23 26 F4 FE 83 27 44 FD
93 97 27 00 23 24 F4 FE 03 27 84 FE 83 27 C4 FE
33 07 F7 00 B7 07 40 03 B3 07 F7 00 23 22 F4 FE
03 27 84 FE 83 27 C4 FE 33 07 F7 00 B7 07 40 03
93 87 07 14 B3 07 F7 00 23 20 F4 FE B7 07 40 00
13 87 C7 39 83 27 C4 FD 93 97 27 00 B3 07 F7 00
83 A7 07 00 13 87 07 00 83 27 44 FE 23 A0 E7 00
B7 07 40 00 13 87 47 3B 83 27 C4 FD 93 97 27 00
B3 07 F7 00 83 A7 07 00 13 87 07 00 83 27 04 FE
23 A0 E7 00 13 00 00 00 03 24 C1 02 13 01 01 03
67 80 00 00 13 01 01 FE 23 2E 81 00 13 04 01 02
23 26 A4 FE 23 24 B4 FE B7 07 C0 00 93 87 07 22
03 27 84 FE 23 A0 E7 00 B7 07 C0 00 93 87 47 23
03 27 C4 FE 23 A0 E7 00 13 00 00 00 03 24 C1 01
13 01 01 02 67 80 00 00 13 01 01 FE 23 2E 81 00
13 04 01 02 23 26 04 FE B7 07 40 03 23 24 F4 FE
23 26 04 FE 6F 00 40 02 83 27 C4 FE 93 97 27 00
03 27 84 FE B3 07 F7 00 23 A0 07 00 83 27 C4 FE
93 87 17 00 23 26 F4 FE 03 27 C4 FE B7 27 00 00
93 87 F7 57 E3 DA E7 FC 13 00 00 00 13 00 00 00
03 24 C1 01 13 01 01 02 67 80 00 00 13 01 01 FC
23 2E 11 02 23 2C 81 02 13 04 01 04 23 26 A4 FC
23 26 04 FE 23 24 04 FE 83 27 C4 FC 63 D6 07 02
83 27 C4 FE 13 87 17 00 23 26 E4 FE 13 07 04 FF
B3 07 F7 00 13 07 D0 02 23 80 E7 FE 83 27 C4 FC
B3 07 F0 40 23 26 F4 FC 83 27 C4 FC 93 05 A0 00
13 85 07 00 EF 00 40 2A 93 07 05 00 13 F7 F7 0F
83 27 C4 FE 93 86 17 00 23 26 D4 FE 13 07 07 03
13 77 F7 0F 93 06 04 FF B3 87 F6 00 23 80 E7 FE
83 27 C4 FC 93 05 A0 00 13 85 07 00 EF 00 80 1E
93 07 05 00 23 26 F4 FC 83 27 C4 FC E3 46 F0 FA
23 24 04 FE 6F 00 00 07 83 27 84 FE 13 07 04 FF
B3 07 F7 00 83 C7 07 FE A3 0F F4 FC 03 27 C4 FE
83 27 84 FE B3 07 F7 40 93 87 F7 FF 13 07 04 FF
B3 07 F7 00 03 C7 07 FE 83 27 84 FE 93 06 04 FF
B3 87 F6 00 23 80 E7 FE 03 27 C4 FE 83 27 84 FE
B3 07 F7 40 93 87 F7 FF 13 07 04 FF B3 07 F7 00
03 47 F4 FD 23 80 E7 FE 83 27 84 FE 93 87 17 00
23 24 F4 FE 83 27 C4 FE 13 D7 F7 01 B3 07 F7 00
93 D7 17 40 13 87 07 00 83 27 84 FE E3 CE E7 F6
B7 07 C0 00 93 87 47 23 83 A7 07 00 23 22 F4 FE
B7 07 C0 00 93 87 07 22 83 A7 07 00 23 20 F4 FE
23 24 04 FE 6F 00 80 06 83 27 84 FE 13 07 04 FF
B3 07 F7 00 83 C7 07 FE 03 26 04 FE 83 25 44 FE
13 85 07 00 EF F0 DF B0 83 27 04 FE 93 87 17 00
23 20 F4 FE 03 27 04 FE 93 07 00 05 63 1A F7 00
23 20 04 FE 83 27 44 FE 93 87 27 00 23 22 F4 FE
03 27 44 FE 93 07 70 07 63 D4 E7 00 23 22 04 FE
83 27 84 FE 93 87 17 00 23 24 F4 FE 03 27 84 FE
83 27 C4 FE E3 4A F7 F8 B7 07 C0 00 93 87 07 22
03 27 04 FE 23 A0 E7 00 B7 07 C0 00 93 87 47 23
03 27 44 FE 23 A0 E7 00 13 00 00 00 83 20 C1 03
03 24 81 03 13 01 01 04 67 80 00 00 13 01 01 FE
23 2E 11 00 23 2C 81 00 13 04 01 02 B7 07 C0 00
83 A7 07 00 23 26 F4 FE 03 27 C4 FE 93 07 40 00
63 1C F7 02 B7 07 40 00 13 85 07 00 EF F0 1F B2
B7 07 40 00 13 85 87 02 EF F0 5F B1 B7 07 40 00
13 85 07 05 EF F0 9F B0 B7 07 40 00 13 85 87 08
EF F0 DF AF 6F 00 80 00 6F 00 00 00 93 07 00 00
13 85 07 00 83 20 C1 01 03 24 81 01 13 01 01 02
67 80 00 00 63 40 05 06 63 C6 05 06 13 86 05 00
93 05 05 00 13 05 F0 FF 63 0C 06 02 93 06 10 00
63 7A B6 00 63 58 C0 00 13 16 16 00 93 96 16 00
E3 6A B6 FE 13 05 00 00 63 E6 C5 00 B3 85 C5 40
33 65 D5 00 93 D6 16 00 13 56 16 00 E3 96 06 FE
67 80 00 00 93 82 00 00 EF F0 5F FB 13 85 05 00
67 80 02 00 33 05 A0 40 63 48 B0 00 B3 05 B0 40
6F F0 DF F9 B3 05 B0 40 93 82 00 00 EF F0 1F F9
33 05 A0 40 67 80 02 00 93 82 00 00 63 CA 05 00
63 4C 05 00 EF F0 9F F7 13 85 05 00 67 80 02 00
B3 05 B0 40 E3 58 05 FE 33 05 A0 40 EF F0 1F F6
33 05 B0 40 67 80 02 00
