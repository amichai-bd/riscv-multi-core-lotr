@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
6F 00 40 0B 67 80 00 00
@00000088
13 01 01 FD 23 26 11 02 23 24 81 02 13 04 01 03
23 2E A4 FC 03 27 C4 FD 93 07 10 00 63 16 F7 00
93 07 10 00 6F 00 00 03 83 27 C4 FD 93 87 F7 FF
13 85 07 00 EF F0 DF FC 93 07 05 00 93 85 07 00
03 25 C4 FD EF 00 80 0B 93 07 05 00 23 26 F4 FE
83 27 C4 FE 13 85 07 00 83 20 C1 02 03 24 81 02
13 01 01 03 67 80 00 00 13 01 01 FE 23 2E 11 00
23 2C 81 00 13 04 01 02 13 05 40 00 EF F0 5F F8
23 26 A4 FE B7 17 40 00 93 87 07 F0 03 27 C4 FE
23 A0 E7 00 13 00 00 00 13 85 07 00 83 20 C1 01
03 24 81 01 13 01 01 02 67 80 00 00 93 00 00 00
13 81 00 00 93 81 00 00 13 82 00 00 93 82 00 00
13 83 00 00 93 83 00 00 13 84 00 00 93 84 00 00
13 85 00 00 93 85 00 00 13 86 00 00 93 86 00 00
13 87 00 00 93 87 00 00 17 11 40 00 13 01 01 D9
13 05 00 00 93 05 00 00 EF F0 1F F7 13 06 05 00
13 05 00 00 93 F6 15 00 63 84 06 00 33 05 C5 00
93 D5 15 00 13 16 16 00 E3 96 05 FE 67 80 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
