@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 40 13 73 00 10 00
@000000A8
13 01 01 FD 23 26 81 02 13 04 01 03 23 2E A4 FC
23 2C B4 FC 83 27 C4 FD 83 A7 07 00 23 26 F4 FE
83 27 84 FD 03 A7 07 00 83 27 C4 FD 23 A0 E7 00
03 27 C4 FE 83 27 84 FD 23 A0 E7 00 13 00 00 00
03 24 C1 02 13 01 01 03 67 80 00 00 13 01 01 FD
23 26 11 02 23 24 81 02 13 04 01 03 23 2E A4 FC
23 2C B4 FC 23 26 04 FE 6F 00 C0 09 23 24 04 FE
6F 00 00 07 83 27 84 FE 93 97 27 00 03 27 C4 FD
B3 07 F7 00 03 A7 07 00 83 27 84 FE 93 87 17 00
93 97 27 00 83 26 C4 FD B3 87 F6 00 83 A7 07 00
63 DA E7 02 83 27 84 FE 93 97 27 00 03 27 C4 FD
B3 06 F7 00 83 27 84 FE 93 87 17 00 93 97 27 00
03 27 C4 FD B3 07 F7 00 93 85 07 00 13 85 06 00
EF F0 1F F3 83 27 84 FE 93 87 17 00 23 24 F4 FE
03 27 84 FD 83 27 C4 FE B3 07 F7 40 93 87 F7 FF
03 27 84 FE E3 40 F7 F8 83 27 C4 FE 93 87 17 00
23 26 F4 FE 83 27 84 FD 93 87 F7 FF 03 27 C4 FE
E3 4E F7 F4 13 00 00 00 13 00 00 00 83 20 C1 02
03 24 81 02 13 01 01 03 67 80 00 00 13 01 01 FB
23 26 11 04 23 24 81 04 13 04 01 05 B7 07 C0 00
83 A7 07 00 23 20 F4 FE 23 26 04 FE 83 27 04 FE
93 87 C7 FF 13 07 70 00 63 6E F7 1C 13 97 27 00
B7 07 40 00 93 87 07 04 B3 07 F7 00 83 A7 07 00
67 80 07 00 13 00 00 00 83 27 C4 FE 13 87 17 00
23 26 E4 FE 13 07 10 03 E3 58 F7 FE B7 17 40 02
93 87 07 90 23 2C F4 FC 93 05 80 00 03 25 84 FD
EF F0 DF EA 13 00 00 00 83 27 C4 FE 13 87 17 00
23 26 E4 FE 13 07 10 03 E3 58 F7 FE 6F 00 80 17
B7 07 40 00 93 87 07 00 83 A8 07 00 03 A8 47 00
03 A5 87 00 83 A5 C7 00 03 A6 07 01 83 A6 47 01
03 A7 87 01 83 A7 C7 01 23 2C 14 FB 23 2E 04 FB
23 20 A4 FC 23 22 B4 FC 23 24 C4 FC 23 26 D4 FC
23 28 E4 FC 23 2A F4 FC 23 24 04 FE 6F 00 C0 03
83 27 84 FE 13 97 27 00 B7 17 40 00 93 87 07 90
33 07 F7 00 83 27 84 FE 93 97 27 00 93 06 04 FF
B3 87 F6 00 83 A7 87 FC 23 20 F7 00 83 27 84 FE
93 87 17 00 23 24 F4 FE 03 27 84 FE 93 07 70 00
E3 D0 E7 FC 6F 00 00 00 6F 00 00 00 6F 00 00 00
B7 07 40 00 93 87 07 02 83 A8 07 00 03 A8 47 00
03 A5 87 00 83 A5 C7 00 03 A6 07 01 83 A6 47 01
03 A7 87 01 83 A7 C7 01 23 2C 14 FB 23 2E 04 FB
23 20 A4 FC 23 22 B4 FC 23 24 C4 FC 23 26 D4 FC
23 28 E4 FC 23 2A F4 FC 23 22 04 FE 6F 00 C0 03
83 27 44 FE 13 97 27 00 B7 17 40 00 93 87 07 90
33 07 F7 00 83 27 44 FE 93 97 27 00 93 06 04 FF
B3 87 F6 00 83 A7 87 FC 23 20 F7 00 83 27 44 FE
93 87 17 00 23 22 F4 FE 03 27 44 FE 93 07 70 00
E3 D0 E7 FC 6F 00 00 00 13 00 00 00 83 27 C4 FE
13 87 17 00 23 26 E4 FE 13 07 10 03 E3 58 F7 FE
B7 17 40 01 93 87 07 90 23 2E F4 FC 93 05 80 00
03 25 C4 FD EF F0 9F D2 6F 00 00 00 6F 00 00 00
6F 00 00 00 93 07 00 00 13 85 07 00 83 20 C1 04
03 24 81 04 13 01 01 05 67 80 00 00
