@00400800
0C 00 00 00 02 00 00 00 00 00 00 00 06 00 00 00
0A 00 00 00 12 00 00 00 64 00 00 00 04 00 00 00
01 00 00 00 02 00 00 00 03 00 00 00 04 00 00 00
05 00 00 00 06 00 00 00 07 00 00 00 08 00 00 00
09 00 00 00 0A 00 00 00 0B 00 00 00 0C 00 00 00
0D 00 00 00 0E 00 00 00 0F 00 00 00 10 00 00 00
0D 00 00 00 0E 00 00 00 0F 00 00 00 10 00 00 00
09 00 00 00 0A 00 00 00 0B 00 00 00 0C 00 00 00
05 00 00 00 06 00 00 00 07 00 00 00 08 00 00 00
01 00 00 00 02 00 00 00 03 00 00 00 04 00 00 00
06 00 00 00 01 00 00 00 00 00 00 00 03 00 00 00
05 00 00 00 09 00 00 00 32 00 00 00 02 00 00 00
98 03 00 00 CC 03 00 00 64 04 00 00 2C 05 00 00
30 05 00 00 C8 05 00 00 FC 05 00 00 4C 06 00 00
