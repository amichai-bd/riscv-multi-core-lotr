@00000000
13 01 01 FE 23 2E 81 00 13 04 01 02 93 07 50 00
23 26 F4 FE 93 07 30 00 23 24 F4 FE 03 27 C4 FE
83 27 84 FE B3 07 F7 02 23 22 F4 FE 93 07 50 00
23 26 F4 FE 93 07 30 00 23 24 F4 FE 03 27 C4 FE
83 27 84 FE B3 07 F7 02 23 22 F4 FE B7 17 00 00
93 87 07 F0 03 27 44 FE 23 A0 E7 00 93 07 00 00
13 85 07 00 03 24 C1 01 13 01 01 02 67 80 00 00
