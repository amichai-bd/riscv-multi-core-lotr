@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
6F 00 00 18 67 80 00 00
@00000088
13 01 01 FC 23 2E 81 02 13 04 01 04 B7 17 40 00
93 87 07 80 83 A5 07 00 03 A6 47 00 83 A6 87 00
03 A7 C7 00 83 A7 07 01 23 26 B4 FC 23 28 C4 FC
23 2A D4 FC 23 2C E4 FC 23 2E F4 FC 23 26 04 FE
23 24 04 FE 93 07 50 00 23 22 F4 FE 23 26 04 FE
6F 00 C0 0C 23 24 04 FE 6F 00 00 0A 83 27 84 FE
93 97 27 00 13 07 04 FF B3 07 F7 00 03 A7 C7 FD
83 27 84 FE 93 87 17 00 93 97 27 00 93 06 04 FF
B3 87 F6 00 83 A7 C7 FD 63 D2 E7 06 83 27 84 FE
93 97 27 00 13 07 04 FF B3 07 F7 00 83 A7 C7 FD
23 20 F4 FE 83 27 84 FE 93 87 17 00 93 97 27 00
13 07 04 FF B3 07 F7 00 03 A7 C7 FD 83 27 84 FE
93 97 27 00 93 06 04 FF B3 87 F6 00 23 AE E7 FC
83 27 84 FE 93 87 17 00 93 97 27 00 13 07 04 FF
B3 07 F7 00 03 27 04 FE 23 AE E7 FC 83 27 84 FE
93 87 17 00 23 24 F4 FE 03 27 44 FE 83 27 C4 FE
B3 07 F7 40 93 87 F7 FF 03 27 84 FE E3 48 F7 F4
83 27 C4 FE 93 87 17 00 23 26 F4 FE 03 27 C4 FE
83 27 44 FE E3 48 F7 F2 B7 17 40 00 03 27 C4 FC
23 A0 E7 00 B7 17 40 00 03 27 04 FD 23 A2 E7 00
B7 17 40 00 03 27 44 FD 23 A4 E7 00 B7 17 40 00
03 27 84 FD 23 A6 E7 00 B7 17 40 00 03 27 C4 FD
23 A8 E7 00 13 00 00 00 13 85 07 00 03 24 C1 03
13 01 01 04 67 80 00 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 17 11 40 00 13 01 41 CC 13 05 00 00
93 05 00 00 EF F0 DF E3 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00
@00400800
01 00 00 00 31 00 00 00 24 00 00 00 32 00 00 00
42 00 00 00
