`define DE10_LITE
`define IMEM_8K
`define DMEM_8K