@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 10 32 73 00 10 00
@000000A8
13 01 01 FE 23 2E 81 00 13 04 01 02 23 26 04 FE
6F 00 00 01 83 27 C4 FE 93 87 17 00 23 26 F4 FE
03 27 C4 FE B7 47 01 00 93 87 F7 87 E3 D4 E7 FE
13 00 00 00 13 00 00 00 03 24 C1 01 13 01 01 02
67 80 00 00 13 01 01 FC 23 2E 81 02 13 04 01 04
23 26 A4 FC 23 24 B4 FC 23 22 C4 FC 83 27 84 FC
93 87 17 14 93 97 17 00 03 27 44 FC B3 07 F7 00
23 22 F4 FE B7 17 00 00 93 87 07 E1 23 20 F4 FE
03 27 C4 FC 93 07 07 00 93 97 27 00 B3 87 E7 00
93 97 47 00 93 87 17 00 23 2E F4 FC 23 26 04 FE
6F 00 40 03 03 27 44 FE 83 27 C4 FE 33 07 F7 40
83 27 04 FE B3 07 F7 00 13 97 27 00 B7 07 40 03
B3 07 F7 00 23 A0 07 00 83 27 C4 FE 93 87 07 05
23 26 F4 FE 03 27 C4 FE B7 17 00 00 93 87 07 96
E3 D2 E7 FC 23 24 04 FE 6F 00 80 03 03 27 44 FE
83 27 84 FE 33 07 F7 40 83 27 04 FE B3 07 F7 00
13 97 27 00 B7 07 40 03 B3 07 F7 00 13 07 F0 FF
23 A0 E7 00 83 27 84 FE 93 87 07 05 23 24 F4 FE
03 27 84 FE 83 27 C4 FD E3 42 F7 FC 13 00 00 00
13 00 00 00 03 24 C1 03 13 01 01 04 67 80 00 00
13 01 01 FD 23 26 81 02 13 04 01 03 23 2E A4 FC
23 2C B4 FC 83 27 C4 FD 83 A7 07 00 23 26 F4 FE
83 27 84 FD 03 A7 07 00 83 27 C4 FD 23 A0 E7 00
83 27 84 FD 03 27 C4 FE 23 A0 E7 00 13 00 00 00
03 24 C1 02 13 01 01 03 67 80 00 00 13 01 01 FD
23 26 11 02 23 24 81 02 13 04 01 03 23 2E A4 FC
23 2C B4 FC 23 2A C4 FC 83 27 44 FD 93 97 27 00
03 27 C4 FD B3 07 F7 00 83 A7 07 00 23 22 F4 FE
83 27 84 FD 93 87 F7 FF 23 26 F4 FE 83 27 84 FD
23 24 F4 FE 6F 00 C0 0D 83 27 84 FE 93 97 27 00
03 27 C4 FD B3 07 F7 00 83 A7 07 00 03 27 44 FE
63 4A F7 0A 83 27 C4 FE 93 87 17 00 23 26 F4 FE
83 27 C4 FE 93 97 27 00 03 27 C4 FD B3 06 F7 00
83 27 84 FE 93 97 27 00 03 27 C4 FD B3 07 F7 00
93 85 07 00 13 85 06 00 EF F0 9F F1 83 27 C4 FE
93 97 27 00 03 27 C4 FD B3 07 F7 00 83 A7 07 00
13 06 40 01 83 25 C4 FE 13 85 07 00 EF F0 9F DF
83 27 84 FE 93 97 27 00 03 27 C4 FD B3 07 F7 00
83 A7 07 00 13 06 40 01 83 25 84 FE 13 85 07 00
EF F0 5F DD 83 27 C4 FE 93 97 27 00 03 27 C4 FD
B3 07 F7 00 03 A7 07 00 83 27 84 FE 93 97 27 00
83 26 C4 FD B3 87 F6 00 83 A7 07 00 63 04 F7 00
EF F0 1F D6 83 27 84 FE 93 87 17 00 23 24 F4 FE
03 27 44 FD 83 27 84 FE E3 C0 E7 F2 83 27 C4 FE
93 87 17 00 93 97 27 00 03 27 C4 FD B3 06 F7 00
83 27 44 FD 93 97 27 00 03 27 C4 FD B3 07 F7 00
93 85 07 00 13 85 06 00 EF F0 9F E5 83 27 C4 FE
93 87 17 00 93 97 27 00 03 27 C4 FD B3 07 F7 00
03 A7 07 00 83 27 C4 FE 93 87 17 00 13 06 40 01
93 85 07 00 13 05 07 00 EF F0 DF D2 83 27 44 FD
93 97 27 00 03 27 C4 FD B3 07 F7 00 83 A7 07 00
13 06 40 01 83 25 44 FD 13 85 07 00 EF F0 9F D0
83 27 C4 FE 93 87 17 00 93 97 27 00 03 27 C4 FD
B3 07 F7 00 03 A7 07 00 83 27 44 FD 93 97 27 00
83 26 C4 FD B3 87 F6 00 83 A7 07 00 63 04 F7 00
EF F0 1F C9 83 27 C4 FE 93 87 17 00 13 85 07 00
83 20 C1 02 03 24 81 02 13 01 01 03 67 80 00 00
13 01 01 FD 23 26 11 02 23 24 81 02 23 22 91 02
13 04 01 03 23 2E A4 FC 23 2C B4 FC 23 2A C4 FC
93 06 01 00 93 84 06 00 03 26 44 FD 83 26 84 FD
B3 06 D6 40 93 86 16 00 13 86 F6 FF 23 24 C4 FE
13 86 06 00 13 0E 06 00 93 0E 00 00 13 56 BE 01
93 98 5E 00 B3 68 16 01 13 18 5E 00 13 86 06 00
13 03 06 00 93 03 00 00 13 56 B3 01 93 97 53 00
B3 67 F6 00 13 17 53 00 93 87 06 00 93 97 27 00
93 87 F7 00 93 D7 47 00 93 97 47 00 33 01 F1 40
93 07 01 00 93 87 37 00 93 D7 27 00 93 97 27 00
23 22 F4 FE 93 07 F0 FF 23 26 F4 FE 83 27 C4 FE
93 87 17 00 23 26 F4 FE 03 27 44 FE 83 27 C4 FE
93 97 27 00 B3 07 F7 00 03 27 84 FD 23 A0 E7 00
83 27 C4 FE 93 87 17 00 23 26 F4 FE 03 27 44 FE
83 27 C4 FE 93 97 27 00 B3 07 F7 00 03 27 44 FD
23 A0 E7 00 6F 00 00 11 83 27 C4 FE 13 87 F7 FF
23 26 E4 FE 03 27 44 FE 93 97 27 00 B3 07 F7 00
83 A7 07 00 23 2A F4 FC 83 27 C4 FE 13 87 F7 FF
23 26 E4 FE 03 27 44 FE 93 97 27 00 B3 07 F7 00
83 A7 07 00 23 2C F4 FC 03 26 44 FD 83 25 84 FD
03 25 C4 FD EF F0 9F CB 23 20 A4 FE 83 27 04 FE
93 87 F7 FF 03 27 84 FD 63 58 F7 04 83 27 C4 FE
93 87 17 00 23 26 F4 FE 03 27 44 FE 83 27 C4 FE
93 97 27 00 B3 07 F7 00 03 27 84 FD 23 A0 E7 00
83 27 C4 FE 93 87 17 00 23 26 F4 FE 83 27 04 FE
13 87 F7 FF 83 26 44 FE 83 27 C4 FE 93 97 27 00
B3 87 F6 00 23 A0 E7 00 83 27 04 FE 93 87 17 00
03 27 44 FD 63 D8 E7 04 83 27 C4 FE 93 87 17 00
23 26 F4 FE 83 27 04 FE 13 87 17 00 83 26 44 FE
83 27 C4 FE 93 97 27 00 B3 87 F6 00 23 A0 E7 00
83 27 C4 FE 93 87 17 00 23 26 F4 FE 03 27 44 FE
83 27 C4 FE 93 97 27 00 B3 07 F7 00 03 27 44 FD
23 A0 E7 00 83 27 C4 FE E3 D8 07 EE 13 81 04 00
13 00 00 00 13 01 04 FD 83 20 C1 02 03 24 81 02
83 24 41 02 13 01 01 03 67 80 00 00 13 01 01 FE
23 2E 81 00 13 04 01 02 23 26 A4 FE 23 24 B4 FE
03 27 C4 FE 83 27 84 FE 63 54 F7 00 93 07 07 00
13 85 07 00 03 24 C1 01 13 01 01 02 67 80 00 00
13 01 01 FD 23 26 11 02 23 24 81 02 13 04 01 03
23 2E A4 FC 23 2C B4 FC 93 07 10 00 23 26 F4 FE
6F 00 40 0A 23 24 04 FE 6F 00 00 08 03 27 84 FE
83 27 C4 FE B3 07 F7 00 13 87 F7 FF 83 27 84 FD
93 87 F7 FF 93 85 07 00 13 05 07 00 EF F0 1F F8
23 22 A4 FE 83 27 C4 FE 13 97 17 00 83 27 84 FE
B3 07 F7 00 13 87 F7 FF 83 27 84 FD 93 87 F7 FF
93 85 07 00 13 05 07 00 EF F0 5F F5 23 20 A4 FE
83 26 04 FE 03 26 44 FE 83 25 84 FE 03 25 C4 FD
EF 00 80 05 83 27 C4 FE 93 97 17 00 03 27 84 FE
B3 07 F7 00 23 24 F4 FE 83 27 84 FD 93 87 F7 FF
03 27 84 FE E3 4C F7 F6 83 27 C4 FE 93 97 17 00
23 26 F4 FE 03 27 84 FD 83 27 C4 FE E3 CC E7 F4
13 00 00 00 13 00 00 00 83 20 C1 02 03 24 81 02
13 01 01 03 67 80 00 00 13 01 01 F9 23 26 11 06
23 24 81 06 23 22 91 06 23 20 21 07 23 2E 31 05
23 2C 41 05 23 2A 51 05 23 28 61 05 23 26 71 05
13 04 01 07 23 2E A4 F8 23 2C B4 F8 23 2A C4 F8
23 28 D4 F8 93 06 01 00 93 84 06 00 03 26 44 F9
83 26 84 F9 B3 06 D6 40 93 86 16 00 23 20 D4 FC
03 26 04 F9 83 26 44 F9 B3 06 D6 40 23 2E D4 FA
83 26 04 FC 13 86 F6 FF 23 2C C4 FA 13 86 06 00
13 0B 06 00 93 0B 00 00 13 56 BB 01 93 9E 5B 00
B3 6E D6 01 13 1E 5B 00 13 86 06 00 13 0A 06 00
93 0A 00 00 13 56 BA 01 93 93 5A 00 B3 63 76 00
13 13 5A 00 93 96 26 00 93 86 F6 00 93 D6 46 00
93 96 46 00 33 01 D1 40 93 06 01 00 93 86 36 00
93 D6 26 00 93 96 26 00 23 2A D4 FA 83 26 C4 FB
13 86 F6 FF 23 28 C4 FA 13 86 06 00 13 09 06 00
93 09 00 00 13 56 B9 01 93 98 59 00 B3 68 16 01
13 18 59 00 13 86 06 00 13 0F 06 00 93 0F 00 00
13 56 BF 01 93 97 5F 00 B3 67 F6 00 13 17 5F 00
93 87 06 00 93 97 27 00 93 87 F7 00 93 D7 47 00
93 97 47 00 33 01 F1 40 93 07 01 00 93 87 37 00
93 D7 27 00 93 97 27 00 23 26 F4 FA 23 22 04 FC
6F 00 00 04 03 27 84 F9 83 27 44 FC B3 07 F7 00
93 97 27 00 03 27 C4 F9 B3 07 F7 00 03 A7 07 00
83 26 44 FB 83 27 44 FC 93 97 27 00 B3 87 F6 00
23 A0 E7 00 83 27 44 FC 93 87 17 00 23 22 F4 FC
03 27 44 FC 83 27 04 FC E3 4E F7 FA 23 24 04 FC
6F 00 40 04 83 27 44 F9 13 87 17 00 83 27 84 FC
B3 07 F7 00 93 97 27 00 03 27 C4 F9 B3 07 F7 00
03 A7 07 00 83 26 C4 FA 83 27 84 FC 93 97 27 00
B3 87 F6 00 23 A0 E7 00 83 27 84 FC 93 87 17 00
23 24 F4 FC 03 27 84 FC 83 27 C4 FB E3 4C F7 FA
23 22 04 FC 23 24 04 FC 83 27 84 F9 23 26 F4 FC
6F 00 00 10 03 27 44 FB 83 27 44 FC 93 97 27 00
B3 07 F7 00 03 A7 07 00 83 26 C4 FA 83 27 84 FC
93 97 27 00 B3 87 F6 00 83 A7 07 00 63 C4 E7 06
83 27 C4 FC 93 97 27 00 03 27 C4 F9 B3 07 F7 00
83 26 44 FB 03 27 44 FC 13 17 27 00 33 87 E6 00
03 27 07 00 23 A0 E7 00 83 27 C4 FC 93 97 27 00
03 27 C4 F9 B3 07 F7 00 03 A7 07 00 B7 17 00 00
13 86 47 2D 83 25 C4 FC 13 05 07 00 EF F0 8F EF
EF F0 0F EB 83 27 44 FC 93 87 17 00 23 22 F4 FC
6F 00 40 06 83 27 C4 FC 93 97 27 00 03 27 C4 F9
B3 07 F7 00 83 26 C4 FA 03 27 84 FC 13 17 27 00
33 87 E6 00 03 27 07 00 23 A0 E7 00 83 27 C4 FC
93 97 27 00 03 27 C4 F9 B3 07 F7 00 03 A7 07 00
B7 17 00 00 13 86 47 2D 83 25 C4 FC 13 05 07 00
EF F0 4F E9 EF F0 CF E4 83 27 84 FC 93 87 17 00
23 24 F4 FC 83 27 C4 FC 93 87 17 00 23 26 F4 FC
03 27 44 FC 83 27 04 FC 63 50 F7 08 03 27 84 FC
83 27 C4 FB E3 48 F7 EE 6F 00 00 07 83 27 C4 FC
93 97 27 00 03 27 C4 F9 B3 07 F7 00 83 26 44 FB
03 27 44 FC 13 17 27 00 33 87 E6 00 03 27 07 00
23 A0 E7 00 83 27 C4 FC 93 97 27 00 03 27 C4 F9
B3 07 F7 00 03 A7 07 00 B7 17 00 00 13 86 47 2D
83 25 C4 FC 13 05 07 00 EF F0 CF E0 EF F0 4F DC
83 27 44 FC 93 87 17 00 23 22 F4 FC 83 27 C4 FC
93 87 17 00 23 26 F4 FC 03 27 44 FC 83 27 04 FC
E3 46 F7 F8 6F 00 00 07 83 27 C4 FC 93 97 27 00
03 27 C4 F9 B3 07 F7 00 83 26 C4 FA 03 27 84 FC
13 17 27 00 33 87 E6 00 03 27 07 00 23 A0 E7 00
83 27 C4 FC 93 97 27 00 03 27 C4 F9 B3 07 F7 00
03 A7 07 00 B7 17 00 00 13 86 47 2D 83 25 C4 FC
13 05 07 00 EF F0 0F D9 EF F0 8F D4 83 27 84 FC
93 87 17 00 23 24 F4 FC 83 27 C4 FC 93 87 17 00
23 26 F4 FC 03 27 84 FC 83 27 C4 FB E3 46 F7 F8
13 81 04 00 13 00 00 00 13 01 04 F9 83 20 C1 06
03 24 81 06 83 24 41 06 03 29 01 06 83 29 C1 05
03 2A 81 05 83 2A 41 05 03 2B 01 05 83 2B C1 04
13 01 01 07 67 80 00 00 13 01 01 F9 23 26 11 06
23 24 81 06 13 04 01 07 B7 07 C0 00 83 A7 07 00
23 20 F4 FE 03 27 04 FE 93 07 70 00 63 08 F7 24
03 27 04 FE 93 07 70 00 63 C8 E7 34 03 27 04 FE
93 07 60 00 63 02 F7 14 03 27 04 FE 93 07 60 00
63 CC E7 32 03 27 04 FE 93 07 40 00 63 0A F7 00
03 27 04 FE 93 07 50 00 63 0E F7 10 6F 00 C0 31
EF F0 0F C8 EF F0 CF C7 EF F0 8F C7 EF F0 4F C7
93 07 B0 00 23 28 F4 F8 93 07 50 00 23 2A F4 F8
93 07 90 00 23 2C F4 F8 93 07 D0 00 23 2E F4 F8
93 07 20 01 23 20 F4 FA 93 07 70 00 23 22 F4 FA
93 07 10 00 23 24 F4 FA 93 07 20 00 23 26 F4 FA
93 07 C0 00 23 28 F4 FA 93 07 A0 00 23 2A F4 FA
93 07 40 00 23 2C F4 FA 93 07 30 00 23 2E F4 FA
93 07 E0 00 23 20 F4 FC 93 07 60 00 23 22 F4 FC
93 07 F0 00 23 24 F4 FC 93 07 10 01 23 26 F4 FC
93 07 80 00 23 28 F4 FC 93 07 00 01 23 2A F4 FC
93 07 20 01 23 2C F4 FC 23 24 04 FE 6F 00 40 03
83 27 84 FE 93 97 27 00 13 07 04 FF B3 07 F7 00
83 A7 07 FA 13 06 40 01 83 25 84 FE 13 85 07 00
EF F0 4F BF 83 27 84 FE 93 87 17 00 23 24 F4 FE
03 27 84 FE 83 27 84 FD E3 44 F7 FC EF F0 4F B9
83 27 84 FD 13 87 F7 FF 93 07 04 F9 13 06 07 00
93 05 00 00 13 85 07 00 EF F0 8F F0 EF F0 4F B7
6F F0 1F EF 6F 00 00 00 23 26 04 FE 6F 00 C0 06
83 27 C4 FE 13 97 27 00 B7 07 40 03 B3 07 F7 00
13 07 F0 FF 23 A0 E7 00 03 27 C4 FE B7 17 00 00
93 87 07 2C B3 07 F7 00 13 97 27 00 B7 07 40 03
93 87 07 EC B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
83 27 C4 FE 13 97 27 00 B7 97 40 03 93 87 07 4C
B3 07 F7 00 13 07 F0 FF 23 A0 E7 00 83 27 C4 FE
93 87 17 00 23 26 F4 FE 03 27 C4 FE 93 07 F0 04
E3 D8 E7 F8 23 26 04 FE 6F 00 40 06 03 27 C4 FE
93 07 07 00 93 97 27 00 B3 87 E7 00 93 97 67 00
13 87 07 00 B7 07 40 03 B3 07 F7 00 13 07 F0 FF
23 A0 E7 00 03 27 C4 FE 93 07 07 00 93 97 27 00
B3 87 E7 00 93 97 67 00 13 87 07 00 B7 07 40 03
93 87 C7 13 B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
83 27 C4 FE 93 87 17 00 23 26 F4 FE 03 27 C4 FE
93 07 70 07 E3 DC E7 F8 6F 00 00 00 EF F0 4F A7
EF F0 0F A7 EF F0 CF A6 EF F0 8F A6 93 07 B0 00
23 28 F4 F8 93 07 50 00 23 2A F4 F8 93 07 90 00
23 2C F4 F8 93 07 D0 00 23 2E F4 F8 93 07 20 01
23 20 F4 FA 93 07 70 00 23 22 F4 FA 93 07 10 00
23 24 F4 FA 93 07 20 00 23 26 F4 FA 93 07 C0 00
23 28 F4 FA 93 07 A0 00 23 2A F4 FA 93 07 40 00
23 2C F4 FA 93 07 30 00 23 2E F4 FA 93 07 E0 00
23 20 F4 FC 93 07 60 00 23 22 F4 FC 93 07 F0 00
23 24 F4 FC 93 07 10 01 23 26 F4 FC 93 07 80 00
23 28 F4 FC 93 07 00 01 23 2A F4 FC 93 07 20 01
23 2E F4 FC 23 22 04 FE 6F 00 80 03 83 27 44 FE
93 97 27 00 13 07 04 FF B3 07 F7 00 03 A7 07 FA
B7 17 00 00 13 86 47 2D 83 25 44 FE 13 05 07 00
EF F0 4F 9E 83 27 44 FE 93 87 17 00 23 22 F4 FE
03 27 44 FE 83 27 C4 FD E3 42 F7 FC EF F0 4F 98
93 07 04 F9 83 25 C4 FD 13 85 07 00 EF F0 4F F6
EF F0 0F 97 6F F0 9F EF 6F 00 00 00
