@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 40 49 73 00 10 00
@000000A8
13 01 01 FE 23 2E 81 00 13 04 01 02 23 26 A4 FE
83 27 C4 FE 93 87 27 0A 13 97 27 00 B7 07 40 03
B3 07 F7 00 13 07 F0 FF 23 A0 E7 00 83 27 C4 FE
93 87 27 0F 13 97 27 00 B7 07 40 03 B3 07 F7 00
13 07 F0 FF 23 A0 E7 00 83 27 C4 FE 93 87 27 14
13 97 27 00 B7 07 40 03 B3 07 F7 00 13 07 F0 FF
23 A0 E7 00 83 27 C4 FE 93 87 27 19 13 97 27 00
B7 07 40 03 B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
83 27 C4 FE 93 87 27 1E 13 97 27 00 B7 07 40 03
B3 07 F7 00 13 07 F0 FF 23 A0 E7 00 83 27 C4 FE
93 87 27 23 13 97 27 00 B7 07 40 03 B3 07 F7 00
13 07 F0 FF 23 A0 E7 00 83 27 C4 FE 93 87 27 28
13 97 27 00 B7 07 40 03 B3 07 F7 00 13 07 F0 FF
23 A0 E7 00 83 27 C4 FE 93 87 47 0A 13 97 27 00
B7 07 40 03 B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
83 27 C4 FE 93 87 47 0F 13 97 27 00 B7 07 40 03
B3 07 F7 00 13 07 F0 FF 23 A0 E7 00 83 27 C4 FE
93 87 47 14 13 97 27 00 B7 07 40 03 B3 07 F7 00
13 07 F0 FF 23 A0 E7 00 83 27 C4 FE 93 87 47 19
13 97 27 00 B7 07 40 03 B3 07 F7 00 13 07 F0 FF
23 A0 E7 00 83 27 C4 FE 93 87 47 1E 13 97 27 00
B7 07 40 03 B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
83 27 C4 FE 93 87 47 23 13 97 27 00 B7 07 40 03
B3 07 F7 00 13 07 F0 FF 23 A0 E7 00 83 27 C4 FE
93 87 47 28 13 97 27 00 B7 07 40 03 B3 07 F7 00
13 07 F0 FF 23 A0 E7 00 83 27 C4 FE 93 87 37 19
13 97 27 00 B7 07 40 03 B3 07 F7 00 13 07 F0 FF
23 A0 E7 00 83 27 C4 FE 93 87 67 0A 13 97 27 00
B7 07 40 03 B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
83 27 C4 FE 93 87 77 0A 13 97 27 00 B7 07 40 03
B3 07 F7 00 13 07 F0 FF 23 A0 E7 00 83 27 C4 FE
93 87 87 0A 13 97 27 00 B7 07 40 03 B3 07 F7 00
13 07 F0 FF 23 A0 E7 00 83 27 C4 FE 93 87 77 0F
13 97 27 00 B7 07 40 03 B3 07 F7 00 13 07 F0 FF
23 A0 E7 00 83 27 C4 FE 93 87 77 14 13 97 27 00
B7 07 40 03 B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
83 27 C4 FE 93 87 77 19 13 97 27 00 B7 07 40 03
B3 07 F7 00 13 07 F0 FF 23 A0 E7 00 83 27 C4 FE
93 87 77 1E 13 97 27 00 B7 07 40 03 B3 07 F7 00
13 07 F0 FF 23 A0 E7 00 83 27 C4 FE 93 87 77 23
13 97 27 00 B7 07 40 03 B3 07 F7 00 13 07 F0 FF
23 A0 E7 00 83 27 C4 FE 93 87 67 28 13 97 27 00
B7 07 40 03 B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
83 27 C4 FE 93 87 77 28 13 97 27 00 B7 07 40 03
B3 07 F7 00 13 07 F0 FF 23 A0 E7 00 83 27 C4 FE
93 87 87 28 13 97 27 00 B7 07 40 03 B3 07 F7 00
13 07 F0 FF 23 A0 E7 00 83 27 C4 FE 93 87 97 19
13 97 27 00 B7 07 40 03 B3 07 F7 00 13 07 F0 FF
23 A0 E7 00 83 27 C4 FE 93 87 A7 19 13 97 27 00
B7 07 40 03 B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
93 07 00 00 13 85 07 00 03 24 C1 01 13 01 01 02
67 80 00 00 13 01 01 FE 23 2E 81 00 13 04 01 02
23 26 A4 FE 83 27 C4 FE 93 87 67 0A 13 97 27 00
B7 07 40 03 B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
83 27 C4 FE 93 87 77 0A 13 97 27 00 B7 07 40 03
B3 07 F7 00 13 07 F0 FF 23 A0 E7 00 83 27 C4 FE
93 87 87 0A 13 97 27 00 B7 07 40 03 B3 07 F7 00
13 07 F0 FF 23 A0 E7 00 83 27 C4 FE 93 87 77 0F
13 97 27 00 B7 07 40 03 B3 07 F7 00 13 07 F0 FF
23 A0 E7 00 83 27 C4 FE 93 87 77 14 13 97 27 00
B7 07 40 03 B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
83 27 C4 FE 93 87 77 19 13 97 27 00 B7 07 40 03
B3 07 F7 00 13 07 F0 FF 23 A0 E7 00 83 27 C4 FE
93 87 77 1E 13 97 27 00 B7 07 40 03 B3 07 F7 00
13 07 F0 FF 23 A0 E7 00 83 27 C4 FE 93 87 77 23
13 97 27 00 B7 07 40 03 B3 07 F7 00 13 07 F0 FF
23 A0 E7 00 83 27 C4 FE 93 87 67 28 13 97 27 00
B7 07 40 03 B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
83 27 C4 FE 93 87 77 28 13 97 27 00 B7 07 40 03
B3 07 F7 00 13 07 F0 FF 23 A0 E7 00 83 27 C4 FE
93 87 87 28 13 97 27 00 B7 07 40 03 B3 07 F7 00
13 07 F0 FF 23 A0 E7 00 93 07 00 00 13 85 07 00
03 24 C1 01 13 01 01 02 67 80 00 00 13 01 01 FE
23 2E 11 00 23 2C 81 00 13 04 01 02 B7 07 C0 00
93 87 47 00 83 A7 07 00 23 24 F4 FE B7 07 C0 00
83 A7 07 00 23 22 F4 FE 23 20 04 FE 03 27 44 FE
93 07 70 00 63 0E F7 1C 03 27 44 FE 93 07 70 00
63 C8 E7 20 03 27 44 FE 93 07 60 00 63 08 F7 18
03 27 44 FE 93 07 60 00 63 CC E7 1E 03 27 44 FE
93 07 40 00 63 0A F7 00 03 27 44 FE 93 07 50 00
63 08 F7 14 6F 00 C0 1D 23 26 04 FE 6F 00 C0 06
83 27 C4 FE 13 97 27 00 B7 07 40 03 B3 07 F7 00
13 07 F0 FF 23 A0 E7 00 03 27 C4 FE B7 17 00 00
93 87 07 2C B3 07 F7 00 13 97 27 00 B7 07 40 03
93 87 07 EC B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
83 27 C4 FE 13 97 27 00 B7 97 40 03 93 87 07 4C
B3 07 F7 00 13 07 F0 FF 23 A0 E7 00 83 27 C4 FE
93 87 17 00 23 26 F4 FE 03 27 C4 FE 93 07 F0 04
E3 D8 E7 F8 23 26 04 FE 6F 00 00 09 03 27 C4 FE
93 07 07 00 93 97 27 00 B3 87 E7 00 93 97 67 00
13 87 07 00 B7 07 40 03 B3 07 F7 00 13 07 F0 FF
23 A0 E7 00 03 27 C4 FE 93 07 07 00 93 97 27 00
B3 87 E7 00 93 97 67 00 13 87 07 00 B7 07 40 03
93 87 C7 09 B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
03 27 C4 FE 93 07 07 00 93 97 27 00 B3 87 E7 00
93 97 67 00 13 87 07 00 B7 07 40 03 93 87 C7 13
B3 07 F7 00 13 07 F0 FF 23 A0 E7 00 83 27 C4 FE
93 87 17 00 23 26 F4 FE 03 27 C4 FE 93 07 70 07
E3 D6 E7 F6 13 05 00 00 EF F0 9F 9D 13 05 60 00
EF F0 5F D0 B7 07 40 03 13 87 47 14 B7 17 40 00
93 87 07 F0 03 27 07 00 23 A0 E7 00 6F 00 80 09
13 05 80 02 EF F0 DF 9A 13 05 E0 02 EF F0 9F CD
13 05 00 03 EF F0 1F CD 6F 00 00 00 B7 17 00 00
13 85 07 2C EF F0 DF 98 B7 17 00 00 13 85 67 2C
EF F0 5F CB B7 17 00 00 13 85 87 2C EF F0 9F CA
B7 17 00 00 13 85 A7 2C EF F0 DF C9 6F 00 00 00
B7 17 00 00 13 85 87 2E EF F0 9F 95 B7 17 00 00
13 85 E7 2E EF F0 1F C8 B7 17 00 00 13 85 07 2F
EF F0 5F C7 B7 17 00 00 13 85 27 2F EF F0 9F C6
B7 17 00 00 13 85 47 2F EF F0 DF C5 6F 00 00 00
6F 00 00 00 93 07 00 00 13 85 07 00 83 20 C1 01
03 24 81 01 13 01 01 02 67 80 00 00
