@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 80 00 73 00 10 00
@000000A8
13 01 01 FA 23 2E 11 04 23 2C 81 04 13 04 01 06
B7 07 40 00 13 87 07 00 93 07 04 FA 93 06 07 00
13 07 00 05 13 06 07 00 93 85 06 00 13 85 07 00
EF 00 C0 02 B7 17 40 00 93 87 07 F0 03 27 04 FE
23 A0 E7 00 93 07 00 00 13 85 07 00 83 20 C1 05
03 24 81 05 13 01 01 06 67 80 00 00 B3 47 B5 00
93 F7 37 00 B3 08 C5 00 63 96 07 06 93 07 30 00
63 F2 C7 06 93 77 35 00 13 07 05 00 63 9A 07 0C
13 F6 C8 FF B3 06 E6 40 93 07 00 02 93 02 00 02
63 C2 D7 06 93 86 05 00 93 07 07 00 63 78 C7 02
03 A8 06 00 93 87 47 00 93 86 46 00 23 AE 07 FF
E3 E8 C7 FE 93 07 F6 FF B3 87 E7 40 93 F7 C7 FF
93 87 47 00 33 07 F7 00 B3 85 F5 00 63 68 17 01
67 80 00 00 13 07 05 00 E3 7C 15 FF 83 C7 05 00
13 07 17 00 93 85 15 00 A3 0F F7 FE E3 68 17 FF
67 80 00 00 83 A6 45 00 83 A7 C5 01 83 AF 05 00
03 AF 85 00 83 AE C5 00 03 AE 05 01 03 A3 45 01
03 A8 85 01 23 22 D7 00 83 A6 05 02 23 20 F7 01
23 24 E7 01 23 26 D7 01 23 28 C7 01 23 2A 67 00
23 2C 07 01 23 2E F7 00 13 07 47 02 B3 07 E6 40
23 2E D7 FE 93 85 45 02 E3 C6 F2 FA 6F F0 9F F4
83 C6 05 00 13 07 17 00 93 77 37 00 A3 0F D7 FE
93 85 15 00 E3 8E 07 F0 83 C6 05 00 13 07 17 00
93 77 37 00 A3 0F D7 FE 93 85 15 00 E3 9A 07 FC
6F F0 1F F0
