@00400000
0C 00 00 00 02 00 00 00 00 00 00 00 06 00 00 00
0A 00 00 00 12 00 00 00 64 00 00 00 04 00 00 00
01 00 00 00 02 00 00 00 03 00 00 00 04 00 00 00
05 00 00 00 06 00 00 00 07 00 00 00 08 00 00 00
09 00 00 00 0A 00 00 00 0B 00 00 00 0C 00 00 00
14 00 00 00 0E 00 00 00 0F 00 00 00 10 00 00 00
0D 00 00 00 0E 00 00 00 0F 00 00 00 10 00 00 00
09 00 00 00 0A 00 00 00 0B 00 00 00 0C 00 00 00
05 00 00 00 06 00 00 00 07 00 00 00 08 00 00 00
01 00 00 00 02 00 00 00 03 00 00 00 04 00 00 00
06 00 00 00 01 00 00 00 00 00 00 00 03 00 00 00
05 00 00 00 09 00 00 00 32 00 00 00 02 00 00 00
50 03 00 00 78 03 00 00 20 04 00 00 F8 04 00 00
FC 04 00 00 A4 05 00 00 CC 05 00 00 10 06 00 00
