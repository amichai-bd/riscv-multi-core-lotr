@00400000
57 45 4C 43 4F 4D 45 20 54 4F 20 54 48 45 20 4C
4F 54 52 20 46 50 47 41 0A 00 00 00 41 20 44 55
41 4C 20 43 4F 52 45 20 38 20 54 48 52 45 41 44
20 46 41 42 52 49 43 20 2E 0A 00 00 50 4C 45 41
53 45 20 55 53 45 20 53 57 49 54 43 48 45 53 20
54 4F 20 53 45 4C 45 43 54 0A 00 00 30 30 31 20
3A 20 53 59 53 54 45 4D 20 49 4E 46 4F 52 4D 41
54 49 4F 4E 0A 00 00 00 30 31 30 20 3A 20 4C 45
44 20 53 48 4F 57 0A 00 31 30 30 20 3A 20 47 52
41 50 48 49 43 20 53 4F 52 54 49 4E 47 0A 00 00
31 30 31 20 3A 20 53 4E 41 4B 45 20 47 41 4D 45
0A 00 00 00 57 45 4C 43 4F 4D 45 20 54 4F 20 54
48 45 20 4C 45 44 20 53 48 4F 57 2E 0A 00 00 00
53 45 54 20 54 48 45 20 46 50 47 41 20 53 57 49
54 43 48 45 53 20 54 4F 20 53 45 4C 45 43 54 20
54 48 45 20 4C 45 44 20 46 55 4E 43 54 49 4F 4E
0A 00 00 00 30 30 30 20 3A 20 41 4C 4C 20 4C 45
44 20 42 4C 49 4E 4B 0A 00 00 00 00 30 30 31 20
3A 20 42 49 4E 41 52 59 20 43 4F 55 4E 54 45 52
20 0A 00 00 30 31 30 20 3A 20 4F 4E 45 20 4C 45
44 20 4D 4F 56 49 4E 47 20 4C 45 46 54 0A 00 00
30 31 31 20 3A 20 44 45 43 52 45 41 53 45 20 42
49 4E 41 52 59 20 43 4F 55 4E 54 45 52 0A 00 00
4C 4F 54 52 20 46 41 42 52 49 43 0A 00 00 00 00
46 50 47 41 20 2E 0A 00 48 57 20 53 59 53 54 45
4D 20 50 52 4F 50 45 52 54 49 45 53 3A 0A 00 00
4E 55 4D 42 45 52 20 4F 46 20 43 4F 52 45 53 3A
20 32 0A 00 4E 55 4D 42 45 52 20 4F 46 20 54 48
52 45 41 44 20 45 41 43 48 20 43 4F 52 45 3A 20
34 0A 00 00 46 50 47 41 20 4D 4F 44 45 4C 20 3A
20 44 45 31 30 4C 49 47 48 54 0A 00 49 4E 53 54
52 55 43 54 49 4F 4E 20 4D 45 4D 4F 52 59 20 53
49 5A 45 20 46 4F 52 20 45 41 43 48 20 43 4F 52
45 20 3A 20 38 20 4B 42 0A 00 00 00 44 41 54 41
20 4D 45 4D 4F 52 59 20 53 49 5A 45 20 46 4F 52
20 45 41 43 48 20 43 4F 52 45 20 3A 20 38 20 4B
42 0A 00 00 56 47 41 20 4D 45 4D 4F 52 59 20 53
49 5A 45 20 3A 20 33 38 20 4B 42 0A 00 00 00 00
53 4F 4D 45 20 43 52 20 46 45 41 54 55 52 45 53
20 3A 20 0A 00 00 00 00 46 52 45 45 5A 45 20 54
48 52 45 41 44 20 50 43 0A 00 00 00 52 45 53 45
54 20 54 48 52 45 41 44 20 50 43 0A 00 00 00 00
43 52 45 41 54 4F 52 53 3A 20 0A 00 41 44 49 20
4C 45 56 59 20 0A 00 00 53 41 41 52 20 4B 41 44
4F 53 48 20 0A 00 00 00 41 4D 49 43 48 41 49 20
42 45 4E 20 44 41 56 49 44 20 0A 00 43 31 20 54
30 2C 20 42 55 42 42 4C 45 20 53 4F 52 54 20 52
41 4E 44 4F 4D 0A 00 00 54 48 45 20 53 4E 41 4B
45 20 47 41 4D 45 20 49 53 20 44 49 53 41 42 4C
45 44 20 44 55 45 20 54 4F 20 4D 45 4D 4F 52 59
20 53 49 5A 45 0A 00 00 43 31 20 54 31 2C 20 42
55 42 42 4C 45 20 53 4F 52 54 20 33 20 55 4E 49
51 55 45 0A 00 00 00 00 43 31 20 54 32 2C 20 42
55 42 42 4C 45 20 53 4F 52 54 20 52 45 56 45 52
53 45 0A 00 43 31 20 54 33 2C 20 42 55 42 42 4C
45 20 53 4F 52 54 20 41 4C 4D 4F 53 54 20 53 4F
52 54 45 44 0A 00 00 00 43 32 20 54 30 20 2C 49
4E 53 45 52 54 49 4F 4E 20 53 4F 52 54 20 52 41
4E 44 4F 4D 0A 00 00 00 43 32 20 54 31 2C 20 49
4E 53 45 52 54 49 4F 4E 20 53 4F 52 54 20 33 20
55 4E 49 51 55 45 0A 00 43 32 20 54 32 2C 20 49
4E 53 45 52 54 49 4F 4E 20 53 4F 52 54 20 52 45
56 45 52 53 45 0A 00 00 43 32 20 54 33 2C 20 49
4E 53 45 52 54 49 4F 4E 20 53 4F 52 54 20 41 4C
4D 4F 53 54 20 53 4F 52 54 45 44 2E 0A 00 00 00
0B 00 00 00 05 00 00 00 09 00 00 00 0D 00 00 00
12 00 00 00 07 00 00 00 01 00 00 00 02 00 00 00
0C 00 00 00 0A 00 00 00 04 00 00 00 03 00 00 00
0E 00 00 00 06 00 00 00 0F 00 00 00 11 00 00 00
08 00 00 00 10 00 00 00 06 00 00 00 12 00 00 00
0C 00 00 00 0C 00 00 00 06 00 00 00 12 00 00 00
12 00 00 00 06 00 00 00 06 00 00 00 0C 00 00 00
0C 00 00 00 12 00 00 00 06 00 00 00 12 00 00 00
06 00 00 00 0C 00 00 00 12 00 00 00 0C 00 00 00
12 00 00 00 11 00 00 00 10 00 00 00 0F 00 00 00
0E 00 00 00 0D 00 00 00 0C 00 00 00 0B 00 00 00
0A 00 00 00 09 00 00 00 08 00 00 00 07 00 00 00
06 00 00 00 05 00 00 00 04 00 00 00 03 00 00 00
02 00 00 00 01 00 00 00 02 00 00 00 03 00 00 00
04 00 00 00 05 00 00 00 06 00 00 00 07 00 00 00
08 00 00 00 09 00 00 00 0A 00 00 00 0B 00 00 00
0C 00 00 00 0D 00 00 00 0E 00 00 00 0F 00 00 00
10 00 00 00 11 00 00 00 12 00 00 00 01 00 00 00
74 0F 00 00 34 10 00 00 74 13 00 00 A0 15 00 00
68 16 00 00 20 17 00 00 E0 17 00 00 98 18 00 00
@00400550
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 3C 62 52 00 18 1C 1A 00 3C 42 40 00 3C 42 40
00 30 28 24 00 7E 02 3E 00 3C 42 02 00 7E 40 30
00 3C 42 42 00 3C 42 42 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 18 3C 66 00 1E 22 3E 00 3C 3E 02
00 1E 3E 22 00 7E 06 06 00 7E 06 06 00 3C 3E 02
00 66 66 66 00 7E 18 18 00 60 60 60 00 46 66 3E
00 06 06 06 00 42 66 5A 00 62 66 6E 00 3C 66 66
00 3E 66 66 00 3C 42 42 00 3E 66 66 00 7C 06 1E
00 7E 18 18 00 66 66 66 00 66 66 66 00 42 42 42
00 66 66 3C 00 66 66 3C 00 7E 20 10 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 18 18 1E 06 00 00 00 00 00 18 18 00
00 00 00 00 4A 46 3C 00 18 18 7E 00 3C 02 7E 00
38 42 3C 00 7E 20 20 00 40 42 3C 00 3E 42 3C 00
08 08 08 00 3C 42 3C 00 7C 40 3E 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 66 7E 66 00 3E 22 1E 00
02 3E 3C 00 22 3E 1E 00 7E 06 7E 00 7E 06 06 00
3A 22 3C 00 7E 66 66 00 18 18 7E 00 66 66 7C 00
3E 66 46 00 06 06 7E 00 5A 42 42 00 76 66 46 00
66 66 3C 00 3E 06 06 00 52 62 7C 00 3E 66 66 00
78 60 3E 00 18 18 18 00 66 7E 3C 00 66 3C 18 00
5A 7E 42 00 3C 66 66 00 18 18 18 00 08 04 7E 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 30 10 38 7C 30 10 38 38
30 10 38 38 30 10 38 7C 30 10 38 38 00 00 00 00
BA 48 84 82 78 AC 48 44 78 28 28 10 BA 38 10 28
7C 38 48 48 00 00 00 00
