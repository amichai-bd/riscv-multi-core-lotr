@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 00 1F
@00000018
13 01 01 FD 23 26 81 02 13 04 01 03 23 2E A4 FC
23 2C B4 FC 83 27 C4 FD 83 A7 07 00 23 26 F4 FE
83 27 84 FD 03 A7 07 00 83 27 C4 FD 23 A0 E7 00
83 27 84 FD 03 27 C4 FE 23 A0 E7 00 13 00 00 00
03 24 C1 02 13 01 01 03 67 80 00 00 13 01 01 FD
23 26 11 02 23 24 81 02 13 04 01 03 23 2E A4 FC
23 2C B4 FC 23 26 04 FE 6F 00 C0 09 23 24 04 FE
6F 00 00 07 83 27 84 FE 93 97 27 00 03 27 C4 FD
B3 07 F7 00 03 A7 07 00 83 27 84 FE 93 87 17 00
93 97 27 00 83 26 C4 FD B3 87 F6 00 83 A7 07 00
63 DA E7 02 83 27 84 FE 93 97 27 00 03 27 C4 FD
B3 06 F7 00 83 27 84 FE 93 87 17 00 93 97 27 00
03 27 C4 FD B3 07 F7 00 93 85 07 00 13 85 06 00
EF F0 1F F3 83 27 84 FE 93 87 17 00 23 24 F4 FE
03 27 84 FD 83 27 C4 FE B3 07 F7 40 93 87 F7 FF
03 27 84 FE E3 40 F7 F8 83 27 C4 FE 93 87 17 00
23 26 F4 FE 83 27 84 FD 93 87 F7 FF 03 27 C4 FE
E3 4E F7 F4 13 00 00 00 13 00 00 00 83 20 C1 02
03 24 81 02 13 01 01 03 67 80 00 00 13 01 01 FC
23 2E 11 02 23 2C 81 02 13 04 01 04 93 07 60 00
23 26 F4 FC 93 07 10 00 23 28 F4 FC 23 2A 04 FC
93 07 30 00 23 2C F4 FC 93 07 50 00 23 2E F4 FC
93 07 90 00 23 20 F4 FE 93 07 20 03 23 22 F4 FE
93 07 20 00 23 24 F4 FE 93 07 C4 FC 93 05 80 00
13 85 07 00 EF F0 9F EC 23 26 04 FE 6F 00 C0 03
83 27 C4 FE 13 97 27 00 B7 17 40 00 93 87 07 F0
33 07 F7 00 83 27 C4 FE 93 97 27 00 93 06 04 FF
B3 87 F6 00 83 A7 C7 FD 23 20 F7 00 83 27 C4 FE
93 87 17 00 23 26 F4 FE 03 27 C4 FE 93 07 70 00
E3 D0 E7 FC 93 07 00 00 13 85 07 00 83 20 C1 03
03 24 81 03 13 01 01 04 67 80 00 00 93 00 00 00
13 81 00 00 93 81 00 00 13 82 00 00 93 82 00 00
13 83 00 00 93 83 00 00 13 84 00 00 93 84 00 00
13 85 00 00 93 85 00 00 13 86 00 00 93 86 00 00
13 87 00 00 93 87 00 00 13 88 00 00 93 88 00 00
13 89 00 00 93 89 00 00 13 8A 00 00 93 8A 00 00
13 8B 00 00 93 8B 00 00 13 8C 00 00 93 8C 00 00
13 8D 00 00 93 8D 00 00 13 8E 00 00 93 8E 00 00
13 8F 00 00 93 8F 00 00 B7 02 C0 00 93 82 C2 00
03 A1 02 00 EF F0 9F EB 73 00 10 00
