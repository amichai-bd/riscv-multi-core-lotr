@00400000
57 45 20 41 52 45 20 54 48 45 20 50 45 4F 50 4C
45 20 54 48 41 54 20 52 55 4C 45 20 54 48 45 20
57 4F 52 4C 44 2E 0A 00 41 20 46 4F 52 43 45 20
52 55 4E 4E 49 4E 47 20 49 4E 20 45 56 45 52 59
20 42 4F 59 20 41 4E 44 20 47 49 52 4C 2E 0A 00
41 4C 4C 20 52 45 4A 4F 49 43 49 4E 47 20 49 4E
20 54 48 45 20 57 4F 52 4C 44 2C 20 54 41 4B 45
20 4D 45 20 4E 4F 57 20 57 45 20 43 41 4E 20 54
52 59 2E 0A 00 00 00 00 30 31 32 33 34 35 36 37
38 39 0A 00 68 04 00 00 C4 04 00 00 DC 04 00 00
F4 04 00 00 0C 05 00 00
@004000A8
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 3C 62 52 00 18 1C 1A 00 3C 42 40 00 3C 42 40
00 30 28 24 00 7E 02 3E 00 3C 42 02 00 7E 40 30
00 3C 42 42 00 3C 42 42 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 18 3C 66 00 1E 22 3E 00 3C 3E 02
00 1E 3E 22 00 7E 06 06 00 7E 06 06 00 3C 3E 02
00 66 66 66 00 7E 18 18 00 60 60 60 00 46 66 3E
00 06 06 06 00 42 66 5A 00 62 66 6E 00 3C 66 66
00 3E 66 66 00 3C 42 42 00 3E 66 66 00 7C 06 1E
00 7E 18 18 00 66 66 66 00 66 66 66 00 42 42 42
00 66 66 3C 00 66 66 3C 00 7E 20 10 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 18 18 1E 06 00 00 00 00 00 18 18 00
00 00 00 00 4A 46 3C 00 18 18 7E 00 3C 02 7E 00
38 42 3C 00 7E 20 20 00 40 42 3C 00 3E 42 3C 00
08 08 08 00 3C 42 3C 00 7C 40 3E 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 66 7E 66 00 3E 22 1E 00
02 3E 3C 00 22 3E 1E 00 7E 06 7E 00 7E 06 06 00
3A 22 3C 00 7E 66 66 00 18 18 7E 00 66 66 7C 00
3E 66 46 00 06 06 7E 00 5A 42 42 00 76 66 46 00
66 66 3C 00 3E 06 06 00 52 62 7C 00 3E 66 66 00
78 60 3E 00 18 18 18 00 66 7E 3C 00 66 3C 18 00
5A 7E 42 00 3C 66 66 00 18 18 18 00 08 04 7E 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 30 10 38 7C 30 10 38 38
30 10 38 38 30 10 38 7C 30 10 38 38 BA 48 84 82
78 AC 48 44 78 28 28 10 BA 38 10 28 7C 38 48 48
