@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 80 00 73 00 10 00
@000000A8
13 01 01 F9 23 26 81 06 13 04 01 07 B7 07 C0 00
83 A7 07 00 23 2C F4 FC 23 26 04 FE 93 07 10 00
23 2A F4 FC 23 24 04 FE 23 22 04 FE 23 20 04 FE
23 2E 04 FC 23 28 04 FC 93 07 00 04 23 28 F4 F8
93 07 90 07 23 2A F4 F8 93 07 40 02 23 2C F4 F8
93 07 00 03 23 2E F4 F8 93 07 90 01 23 20 F4 FA
93 07 20 01 23 22 F4 FA 93 07 20 00 23 24 F4 FA
93 07 80 07 23 26 F4 FA 23 28 04 FA 93 07 80 01
23 2A F4 FA 93 07 80 00 23 2C F4 FA 93 07 30 00
23 2E F4 FA 93 07 60 04 23 20 F4 FC 93 07 10 02
23 22 F4 FC 93 07 60 00 23 24 F4 FC 93 07 E0 00
23 26 F4 FC 93 07 F0 07 23 28 F4 FC 03 27 84 FD
93 07 70 00 63 0C F7 14 03 27 84 FD 93 07 70 00
63 CC E7 18 03 27 84 FD 93 07 60 00 63 04 F7 0E
03 27 84 FD 93 07 60 00 63 C0 E7 18 03 27 84 FD
93 07 40 00 63 0C F7 06 03 27 84 FD 93 07 50 00
63 14 F7 16 6F 00 00 01 83 27 C4 FE 93 87 17 00
23 26 F4 FE 03 27 C4 FE 93 07 90 0F E3 D6 E7 FE
83 27 84 FE 13 87 17 00 23 24 E4 FE 37 27 C0 03
13 07 07 01 93 97 27 00 93 87 07 FF B3 87 87 00
83 A7 07 FA 23 20 F7 00 03 27 84 FE 93 07 00 01
63 D4 E7 00 23 24 04 FE 23 26 04 FE 6F F0 9F FB
83 27 C4 FE 93 87 17 00 23 26 F4 FE 03 27 C4 FE
93 07 90 0F E3 D6 E7 FE 83 27 44 FE 13 87 17 00
23 22 E4 FE 37 27 C0 03 13 07 47 00 93 97 27 00
93 87 07 FF B3 87 87 00 83 A7 07 FA 23 20 F7 00
03 27 44 FE 93 07 00 01 63 D4 E7 00 23 22 04 FE
23 26 04 FE 6F F0 9F FB 83 27 C4 FE 93 87 17 00
23 26 F4 FE 03 27 C4 FE 93 07 90 0F E3 D6 E7 FE
83 27 04 FE 13 87 17 00 23 20 E4 FE 37 27 C0 03
13 07 87 00 93 97 27 00 93 87 07 FF B3 87 87 00
83 A7 07 FA 23 20 F7 00 03 27 04 FE 93 07 00 01
63 D4 E7 00 23 20 04 FE 23 26 04 FE 6F F0 9F FB
83 27 C4 FE 93 87 17 00 23 26 F4 FE 03 27 C4 FE
93 07 90 0F E3 D6 E7 FE 83 27 C4 FD 13 87 17 00
23 2E E4 FC 37 27 C0 03 13 07 C7 00 93 97 27 00
93 87 07 FF B3 87 87 00 83 A7 07 FA 23 20 F7 00
03 27 C4 FD 93 07 00 01 63 D4 E7 00 23 2E 04 FC
23 26 04 FE 6F F0 9F FB 6F 00 00 00
