@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 10 C0 37 73 00 10 00
@000000A8
13 01 01 FD 23 26 81 02 13 04 01 03 93 07 05 00
23 2C B4 FC 23 2A C4 FC A3 0F F4 FC 03 27 84 FD
93 07 07 00 93 97 27 00 B3 87 E7 00 93 97 67 00
23 26 F4 FE 83 27 44 FD 93 97 27 00 23 24 F4 FE
03 27 84 FE 83 27 C4 FE 33 07 F7 00 B7 07 40 03
B3 07 F7 00 23 22 F4 FE 03 27 84 FE 83 27 C4 FE
33 07 F7 00 B7 07 40 03 93 87 07 14 B3 07 F7 00
23 20 F4 FE 83 47 F4 FD 37 07 40 00 13 07 C7 52
93 97 27 00 B3 07 F7 00 83 A7 07 00 13 87 07 00
83 27 44 FE 23 A0 E7 00 83 47 F4 FD 37 07 40 00
13 07 07 6B 93 97 27 00 B3 07 F7 00 83 A7 07 00
13 87 07 00 83 27 04 FE 23 A0 E7 00 13 00 00 00
03 24 C1 02 13 01 01 03 67 80 00 00 13 01 01 FD
23 26 11 02 23 24 81 02 13 04 01 03 23 2E A4 FC
23 26 04 FE 23 24 04 FE 23 22 04 FE B7 07 C0 00
93 87 07 22 83 A7 07 00 23 22 F4 FE B7 07 C0 00
93 87 47 23 83 A7 07 00 23 24 F4 FE 6F 00 80 0B
83 27 C4 FE 03 27 C4 FD B3 07 F7 00 03 C7 07 00
93 07 A0 00 63 1A F7 02 23 22 04 FE 83 27 84 FE
93 87 27 00 23 24 F4 FE 03 27 84 FE 93 07 80 07
63 14 F7 00 23 24 04 FE 83 27 C4 FE 93 87 17 00
23 26 F4 FE 6F 00 00 07 83 27 C4 FE 03 27 C4 FD
B3 07 F7 00 83 C7 07 00 03 27 84 FE 83 26 44 FE
13 86 06 00 93 05 07 00 13 85 07 00 EF F0 5F E8
83 27 44 FE 93 87 17 00 23 22 F4 FE 03 27 44 FE
93 07 00 05 63 12 F7 02 23 22 04 FE 83 27 84 FE
93 87 27 00 23 24 F4 FE 03 27 84 FE 93 07 80 07
63 14 F7 00 23 24 04 FE 83 27 C4 FE 93 87 17 00
23 26 F4 FE 83 27 C4 FE 03 27 C4 FD B3 07 F7 00
83 C7 07 00 E3 9E 07 F2 B7 07 C0 00 93 87 07 22
03 27 44 FE 23 A0 E7 00 B7 07 C0 00 93 87 47 23
03 27 84 FE 23 A0 E7 00 13 00 00 00 83 20 C1 02
03 24 81 02 13 01 01 03 67 80 00 00 13 01 01 FD
23 26 81 02 13 04 01 03 23 2E A4 FC 23 2C B4 FC
23 2A C4 FC 03 27 84 FD 93 07 07 00 93 97 27 00
B3 87 E7 00 93 97 67 00 23 26 F4 FE 83 27 44 FD
93 97 27 00 23 24 F4 FE 03 27 84 FE 83 27 C4 FE
33 07 F7 00 B7 07 40 03 B3 07 F7 00 23 22 F4 FE
03 27 84 FE 83 27 C4 FE 33 07 F7 00 B7 07 40 03
93 87 07 14 B3 07 F7 00 23 20 F4 FE B7 17 40 00
13 87 47 83 83 27 C4 FD 93 97 27 00 B3 07 F7 00
83 A7 07 00 13 87 07 00 83 27 44 FE 23 A0 E7 00
B7 17 40 00 13 87 C7 84 83 27 C4 FD 93 97 27 00
B3 07 F7 00 83 A7 07 00 13 87 07 00 83 27 04 FE
23 A0 E7 00 13 00 00 00 03 24 C1 02 13 01 01 03
67 80 00 00 13 01 01 FE 23 2E 81 00 13 04 01 02
23 26 A4 FE 23 24 B4 FE B7 07 C0 00 93 87 07 22
03 27 84 FE 23 A0 E7 00 B7 07 C0 00 93 87 47 23
03 27 C4 FE 23 A0 E7 00 13 00 00 00 03 24 C1 01
13 01 01 02 67 80 00 00 13 01 01 FE 23 2E 81 00
13 04 01 02 23 26 04 FE B7 07 40 03 23 24 F4 FE
23 26 04 FE 6F 00 40 02 83 27 C4 FE 93 97 27 00
03 27 84 FE B3 07 F7 00 23 A0 07 00 83 27 C4 FE
93 87 17 00 23 26 F4 FE 03 27 C4 FE B7 27 00 00
93 87 F7 57 E3 DA E7 FC 13 00 00 00 13 00 00 00
03 24 C1 01 13 01 01 02 67 80 00 00 13 01 01 FE
23 2E 81 00 13 04 01 02 23 26 04 FE 6F 00 00 01
83 27 C4 FE 93 87 17 00 23 26 F4 FE 03 27 C4 FE
B7 47 01 00 93 87 F7 87 E3 D4 E7 FE 13 00 00 00
13 00 00 00 03 24 C1 01 13 01 01 02 67 80 00 00
13 01 01 FD 23 26 81 02 13 04 01 03 23 2E A4 FC
23 2C B4 FC 23 2A C4 FC 23 28 D4 FC 83 27 84 FD
93 87 17 14 93 97 17 00 03 27 44 FD B3 07 F7 00
23 22 F4 FE 03 27 C4 FD 93 07 07 00 93 97 27 00
B3 87 E7 00 93 97 47 00 93 87 17 00 23 20 F4 FE
23 26 04 FE 6F 00 40 03 03 27 44 FE 83 27 C4 FE
33 07 F7 40 83 27 04 FD B3 07 F7 00 13 97 27 00
B7 07 40 03 B3 07 F7 00 23 A0 07 00 83 27 C4 FE
93 87 07 05 23 26 F4 FE 03 27 C4 FE 93 07 00 64
E3 D4 E7 FC 23 24 04 FE 6F 00 80 03 03 27 44 FE
83 27 84 FE 33 07 F7 40 83 27 04 FD B3 07 F7 00
13 97 27 00 B7 07 40 03 B3 07 F7 00 13 07 F0 FF
23 A0 E7 00 83 27 84 FE 93 87 07 05 23 24 F4 FE
03 27 84 FE 83 27 04 FE E3 42 F7 FC 13 00 00 00
13 00 00 00 03 24 C1 02 13 01 01 03 67 80 00 00
13 01 01 FD 23 26 81 02 13 04 01 03 23 2E A4 FC
23 2C B4 FC 83 27 C4 FD 83 A7 07 00 23 26 F4 FE
83 27 84 FD 03 A7 07 00 83 27 C4 FD 23 A0 E7 00
83 27 84 FD 03 27 C4 FE 23 A0 E7 00 13 00 00 00
03 24 C1 02 13 01 01 03 67 80 00 00 13 01 01 FD
23 26 11 02 23 24 81 02 13 04 01 03 23 2E A4 FC
23 2C B4 FC 23 2A C4 FC 23 28 D4 FC 23 26 04 FE
6F 00 C0 0F 23 24 04 FE 6F 00 00 0D 83 27 84 FE
93 97 27 00 03 27 C4 FD B3 07 F7 00 03 A7 07 00
83 27 84 FE 93 87 17 00 93 97 27 00 83 26 C4 FD
B3 87 F6 00 83 A7 07 00 63 DA E7 08 83 27 84 FE
93 97 27 00 03 27 C4 FD B3 06 F7 00 83 27 84 FE
93 87 17 00 93 97 27 00 03 27 C4 FD B3 07 F7 00
93 85 07 00 13 85 06 00 EF F0 9F F2 83 27 84 FE
93 97 27 00 03 27 C4 FD B3 07 F7 00 83 A7 07 00
83 26 04 FD 03 26 44 FD 83 25 84 FE 13 85 07 00
EF F0 1F E1 83 27 84 FE 93 87 17 00 93 97 27 00
03 27 C4 FD B3 07 F7 00 03 A7 07 00 83 27 84 FE
93 87 17 00 83 26 04 FD 03 26 44 FD 93 85 07 00
13 05 07 00 EF F0 DF DD EF F0 5F D9 83 27 84 FE
93 87 17 00 23 24 F4 FE 03 27 84 FD 83 27 C4 FE
B3 07 F7 40 93 87 F7 FF 03 27 84 FE E3 40 F7 F2
83 27 C4 FE 93 87 17 00 23 26 F4 FE 83 27 84 FD
93 87 F7 FF 03 27 C4 FE E3 4E F7 EE 13 00 00 00
13 00 00 00 83 20 C1 02 03 24 81 02 13 01 01 03
67 80 00 00 13 01 01 FD 23 26 11 02 23 24 81 02
13 04 01 03 23 2E A4 FC 23 2C B4 FC 23 2A C4 FC
23 28 D4 FC 93 07 10 00 23 26 F4 FE 6F 00 00 12
83 27 C4 FE 93 97 27 00 03 27 C4 FD B3 07 F7 00
83 A7 07 00 23 22 F4 FE 83 27 C4 FE 93 87 F7 FF
23 24 F4 FE 6F 00 40 07 83 27 84 FE 93 97 27 00
03 27 C4 FD 33 07 F7 00 83 27 84 FE 93 87 17 00
93 97 27 00 83 26 C4 FD B3 87 F6 00 03 27 07 00
23 A0 E7 00 83 27 84 FE 93 87 17 00 93 97 27 00
03 27 C4 FD B3 07 F7 00 03 A7 07 00 83 27 84 FE
93 87 17 00 83 26 04 FD 03 26 44 FD 93 85 07 00
13 05 07 00 EF F0 DF CC EF F0 5F C8 83 27 84 FE
93 87 F7 FF 23 24 F4 FE 83 27 84 FE 63 C0 07 02
83 27 84 FE 93 97 27 00 03 27 C4 FD B3 07 F7 00
83 A7 07 00 03 27 44 FE E3 48 F7 F6 83 27 84 FE
93 87 17 00 93 97 27 00 03 27 C4 FD B3 07 F7 00
03 27 44 FE 23 A0 E7 00 83 27 84 FE 93 87 17 00
93 97 27 00 03 27 C4 FD B3 07 F7 00 03 A7 07 00
83 27 84 FE 93 87 17 00 83 26 04 FD 03 26 44 FD
93 85 07 00 13 05 07 00 EF F0 9F C4 EF F0 1F C0
83 27 C4 FE 93 87 17 00 23 26 F4 FE 03 27 C4 FE
83 27 84 FD E3 4E F7 EC 13 00 00 00 13 00 00 00
83 20 C1 02 03 24 81 02 13 01 01 03 67 80 00 00
13 01 01 FF 23 26 11 00 23 24 81 00 13 04 01 01
93 05 10 00 13 05 10 00 EF F0 DF B0 B7 07 40 00
13 85 07 00 EF F0 9F 8F 93 05 10 00 13 05 A0 00
EF F0 5F AF B7 07 40 00 13 85 C7 01 EF F0 1F 8E
93 05 40 01 13 05 40 01 EF F0 DF AD B7 07 40 00
13 85 C7 03 EF F0 9F 8C 93 05 40 01 13 05 80 02
EF F0 5F AC B7 07 40 00 13 85 C7 05 EF F0 1F 8B
93 05 40 01 13 05 20 03 EF F0 DF AA B7 07 40 00
13 85 87 07 EF F0 9F 89 93 05 40 01 13 05 C0 03
EF F0 5F A9 B7 07 40 00 13 85 87 08 EF F0 1F 88
93 05 40 01 13 05 60 04 EF F0 DF A7 B7 07 40 00
13 85 07 0A EF F0 9F 86 13 00 00 00 83 20 C1 00
03 24 81 00 13 01 01 01 67 80 00 00 13 01 01 FD
23 26 11 02 23 24 81 02 13 04 01 03 93 07 10 00
23 26 F4 FE 93 07 F0 3F 23 24 F4 FE 23 22 04 FE
93 07 10 00 23 20 F4 FE 93 07 00 20 23 2E F4 FC
93 05 A0 00 13 05 40 01 EF F0 DF A1 B7 07 40 00
13 85 47 0B EF F0 9F 80 93 05 F0 00 13 05 E0 01
EF F0 5F A0 B7 07 40 00 13 85 07 0D EF F0 0F FF
93 05 40 01 13 05 80 02 EF F0 DF 9E B7 07 40 00
13 85 47 10 EF F0 8F FD 93 05 40 01 13 05 D0 02
EF F0 5F 9D B7 07 40 00 13 85 C7 11 EF F0 0F FC
93 05 40 01 13 05 20 03 EF F0 DF 9B B7 07 40 00
13 85 47 13 EF F0 8F FA 93 05 40 01 13 05 70 03
EF F0 5F 9A B7 07 40 00 13 85 07 15 EF F0 0F F9
B7 27 C0 03 93 87 47 02 83 A7 07 00 63 9C 07 04
93 07 10 00 23 26 F4 FE 93 07 F0 3F 23 24 F4 FE
93 07 10 00 23 20 F4 FE 93 07 00 20 23 2E F4 FC
EF F0 DF A0 B7 27 C0 03 93 87 87 01 03 27 44 FE
23 A0 E7 00 03 27 44 FE 93 07 F0 3F 63 16 F7 00
23 22 04 FE 6F F0 DF FA 93 07 F0 3F 23 22 F4 FE
6F F0 1F FA B7 27 C0 03 93 87 47 02 03 A7 07 00
93 07 10 00 63 1C F7 04 93 07 F0 3F 23 24 F4 FE
23 22 04 FE 93 07 10 00 23 20 F4 FE 93 07 00 20
23 2E F4 FC EF F0 9F 9A B7 27 C0 03 93 87 87 01
03 27 C4 FE 23 A0 E7 00 83 27 C4 FE 93 87 17 00
23 26 F4 FE 03 27 C4 FE 93 07 F0 3F E3 12 F7 F4
93 07 10 00 23 26 F4 FE 6F F0 9F F3 B7 27 C0 03
93 87 47 02 03 A7 07 00 93 07 20 00 63 1C F7 04
93 07 10 00 23 26 F4 FE 93 07 F0 3F 23 24 F4 FE
23 22 04 FE 93 07 00 20 23 2E F4 FC EF F0 1F 94
B7 27 C0 03 93 87 87 01 03 27 04 FE 23 A0 E7 00
83 27 04 FE 93 97 17 00 23 20 F4 FE 03 27 04 FE
93 07 00 20 E3 DE E7 EC 93 07 10 00 23 20 F4 FE
6F F0 1F ED B7 27 C0 03 93 87 47 02 03 A7 07 00
93 07 30 00 E3 1E F7 EA 93 07 10 00 23 26 F4 FE
23 22 04 FE 93 07 10 00 23 20 F4 FE 93 07 00 20
23 2E F4 FC EF F0 9F 8D B7 27 C0 03 93 87 87 01
03 27 84 FE 23 A0 E7 00 83 27 84 FE 93 87 F7 FF
23 24 F4 FE 83 27 84 FE E3 9C 07 E6 93 07 F0 3F
23 24 F4 FE 6F F0 DF E6 13 01 01 FF 23 26 11 00
23 24 81 00 13 04 01 01 93 05 10 00 13 05 10 00
EF F0 4F FE B7 07 40 00 13 85 07 17 EF F0 0F DD
93 05 10 00 13 05 50 00 EF F0 CF FC B7 07 40 00
13 85 07 18 EF F0 8F DB 93 05 40 01 13 05 A0 00
EF F0 4F FB B7 07 40 00 13 85 87 18 EF F0 0F DA
93 05 40 01 13 05 40 01 EF F0 CF F9 B7 07 40 00
13 85 07 1A EF F0 8F D8 93 05 40 01 13 05 90 01
EF F0 4F F8 B7 07 40 00 13 85 47 1B EF F0 0F D7
93 05 40 01 13 05 E0 01 EF F0 CF F6 B7 07 40 00
13 85 47 1D EF F0 8F D5 93 05 40 01 13 05 30 02
EF F0 4F F5 B7 07 40 00 13 85 C7 1E EF F0 0F D4
93 05 40 01 13 05 80 02 EF F0 CF F3 B7 07 40 00
13 85 C7 21 EF F0 8F D2 93 05 40 01 13 05 D0 02
EF F0 4F F2 B7 07 40 00 13 85 47 24 EF F0 0F D1
93 05 40 01 13 05 20 03 EF F0 CF F0 B7 07 40 00
13 85 07 26 EF F0 8F CF 93 05 90 01 13 05 70 03
EF F0 4F EF B7 07 40 00 13 85 87 27 EF F0 0F CE
93 05 90 01 13 05 C0 03 EF F0 CF ED B7 07 40 00
13 85 C7 28 EF F0 8F CC 93 05 40 01 13 05 10 04
EF F0 4F EC B7 07 40 00 13 85 07 2A EF F0 0F CB
93 05 90 01 13 05 60 04 EF F0 CF EA B7 07 40 00
13 85 C7 2A EF F0 8F C9 93 05 90 01 13 05 B0 04
EF F0 4F E9 B7 07 40 00 13 85 87 2B EF F0 0F C8
93 05 90 01 13 05 00 05 EF F0 CF E7 B7 07 40 00
13 85 87 2C EF F0 8F C6 13 00 00 00 83 20 C1 00
03 24 81 00 13 01 01 01 67 80 00 00 13 01 01 FD
23 26 81 02 13 04 01 03 93 07 05 00 A3 0F F4 FC
B7 27 C0 03 93 87 47 02 83 A7 07 00 A3 07 F4 FE
83 47 F4 FE 63 84 07 02 03 47 F4 FE 93 07 20 00
63 0E F7 00 03 47 F4 FE 93 07 40 00 63 08 F7 00
03 47 F4 FE 93 07 10 00 63 1E F7 04 83 47 F4 FD
63 98 07 00 03 47 F4 FE 93 07 40 00 63 04 F7 04
03 47 F4 FD 93 07 40 00 63 16 F7 00 83 47 F4 FE
63 8A 07 02 03 47 F4 FD 93 07 20 00 63 18 F7 00
03 47 F4 FE 93 07 10 00 63 0E F7 00 03 47 F4 FD
93 07 10 00 63 1C F7 00 03 47 F4 FE 93 07 20 00
63 16 F7 00 83 47 F4 FD A3 07 F4 FE 83 47 F4 FE
13 85 07 00 03 24 C1 02 13 01 01 03 67 80 00 00
13 01 01 FD 23 26 81 02 13 04 01 03 93 07 05 00
23 2C B4 FC 23 2A C4 FC 13 87 06 00 A3 0F F4 FC
93 07 07 00 23 0F F4 FC 83 47 E4 FD 93 87 F7 FF
23 26 F4 FE 6F 00 80 05 83 27 C4 FE 93 87 F7 FF
03 27 84 FD 33 07 F7 00 83 27 C4 FE 83 26 84 FD
B3 87 F6 00 03 47 07 00 23 80 E7 00 83 27 C4 FE
93 87 F7 FF 03 27 44 FD 33 07 F7 00 83 27 C4 FE
83 26 44 FD B3 87 F6 00 03 47 07 00 23 80 E7 00
83 27 C4 FE 93 87 F7 FF 23 26 F4 FE 83 27 C4 FE
E3 44 F0 FA 03 47 F4 FD 93 07 20 00 63 18 F7 02
83 27 84 FD 03 C7 17 00 83 27 84 FD 23 80 E7 00
83 27 44 FD 93 87 17 00 83 C7 07 00 93 87 F7 FF
13 F7 F7 0F 83 27 44 FD 23 80 E7 00 03 47 F4 FD
93 07 10 00 63 18 F7 02 83 27 84 FD 03 C7 17 00
83 27 84 FD 23 80 E7 00 83 27 44 FD 93 87 17 00
83 C7 07 00 93 87 17 00 13 F7 F7 0F 83 27 44 FD
23 80 E7 00 03 47 F4 FD 93 07 40 00 63 18 F7 02
83 27 84 FD 93 87 17 00 83 C7 07 00 93 87 F7 FF
13 F7 F7 0F 83 27 84 FD 23 80 E7 00 83 27 44 FD
03 C7 17 00 83 27 44 FD 23 80 E7 00 83 47 F4 FD
63 98 07 02 83 27 84 FD 93 87 17 00 83 C7 07 00
93 87 17 00 13 F7 F7 0F 83 27 84 FD 23 80 E7 00
83 27 44 FD 03 C7 17 00 83 27 44 FD 23 80 E7 00
83 47 F4 FD 63 98 07 02 83 27 84 FD 93 87 17 00
83 C7 07 00 93 87 17 00 13 F7 F7 0F 83 27 84 FD
23 80 E7 00 83 27 44 FD 03 C7 17 00 83 27 44 FD
23 80 E7 00 13 00 00 00 03 24 C1 02 13 01 01 03
67 80 00 00 13 01 01 FD 23 26 11 02 23 24 81 02
13 04 01 03 93 07 05 00 23 2C B4 FC 23 2A C4 FC
23 28 D4 FC A3 0F F4 FC 93 07 07 00 23 0F F4 FC
23 26 04 FE 6F 00 40 0D 83 27 C4 FE 03 27 84 FD
B3 07 F7 00 83 C7 07 00 63 8A 07 0A 83 27 C4 FE
03 27 04 FD B3 07 F7 00 83 C7 07 00 93 96 17 00
83 27 C4 FE 03 27 44 FD B3 07 F7 00 83 C7 07 00
13 86 07 00 93 85 06 00 13 05 80 05 EF F0 4F 89
83 27 C4 FE 93 87 17 00 03 27 84 FD B3 07 F7 00
83 C7 07 00 63 94 07 06 83 47 F4 FD 63 82 07 02
83 27 C4 FE 93 87 17 00 03 27 84 FD B3 07 F7 00
13 07 10 00 23 80 E7 00 A3 0F 04 FC 6F 00 00 04
83 27 C4 FE 93 87 17 00 03 27 04 FD B3 07 F7 00
83 C7 07 00 93 96 17 00 83 27 C4 FE 93 87 17 00
03 27 44 FD B3 07 F7 00 83 C7 07 00 13 86 07 00
93 85 06 00 13 05 00 02 EF F0 8F 81 83 27 C4 FE
93 87 17 00 23 26 F4 FE 83 47 E4 FD 03 27 C4 FE
E3 44 F7 F2 13 00 00 00 13 00 00 00 83 20 C1 02
03 24 81 02 13 01 01 03 67 80 00 00 13 01 01 FD
23 26 81 02 13 04 01 03 23 2E A4 FC 23 2A F4 FC
93 87 05 00 A3 0D F4 FC 93 07 06 00 23 0D F4 FC
93 87 06 00 A3 0C F4 FC 93 07 07 00 23 0C F4 FC
03 47 B4 FD 83 47 94 FD 63 1C F7 00 03 47 A4 FD
83 47 84 FD 63 16 F7 00 93 07 10 00 6F 00 80 00
93 07 00 00 A3 07 F4 FE 83 47 F4 FE 63 8E 07 00
83 27 44 FD 83 C7 07 00 93 87 17 00 13 F7 F7 0F
83 27 44 FD 23 80 E7 00 83 47 F4 FE 13 85 07 00
03 24 C1 02 13 01 01 03 67 80 00 00 13 01 01 FA
23 2E 11 04 23 2C 81 04 13 04 01 06 A3 07 04 FE
93 07 50 00 23 07 F4 FE 93 07 50 00 A3 06 F4 FE
A3 05 04 FA 23 06 04 FE A3 05 04 FE 23 05 04 FE
B7 27 C0 03 93 87 47 02 83 A7 07 00 23 0F F4 FC
83 07 E4 FD 63 D2 07 12 EF F0 0F A2 93 07 50 00
23 07 F4 FE 93 07 50 00 A3 06 F4 FE A3 05 04 FA
23 06 04 FE A3 05 04 FE 23 05 04 FE 23 22 04 FE
6F 00 00 03 03 26 44 FE 93 05 00 00 13 05 10 04
EF E0 1F ED 03 26 44 FE 93 05 60 07 13 05 10 04
EF E0 1F EC 83 27 44 FE 93 87 17 00 23 22 F4 FE
03 27 44 FE 93 07 F0 04 E3 D6 E7 FC 23 20 04 FE
6F 00 00 04 83 27 04 FE 93 97 17 00 13 06 00 00
93 85 07 00 13 05 10 04 EF E0 9F E8 83 27 04 FE
93 97 17 00 13 06 F0 04 93 85 07 00 13 05 10 04
EF E0 1F E7 83 27 04 FE 93 87 17 00 23 20 F4 FE
03 27 04 FE 93 07 B0 03 E3 DE E7 FA A3 0F 04 FC
6F 00 C0 05 83 47 F4 FD 03 47 F4 FD 13 07 47 01
13 77 F7 0F 93 06 04 FF B3 87 F6 00 23 8E E7 FC
83 47 F4 FD 13 07 04 FF B3 07 F7 00 13 07 40 01
23 86 E7 FC 83 47 F4 FD 93 B7 57 00 13 F7 F7 0F
83 47 F4 FD 93 06 04 FF B3 87 F6 00 23 8E E7 FA
83 47 F4 FD 93 87 17 00 A3 0F F4 FC 03 47 F4 FD
93 07 E0 00 E3 F0 E7 FA 83 47 F4 FE 13 85 07 00
EF F0 DF A5 93 07 05 00 A3 07 F4 FE 83 47 B4 FE
63 90 07 02 13 06 C4 FB 13 07 C4 FC 83 47 F4 FE
93 06 F0 00 93 05 07 00 13 85 07 00 EF F0 5F AF
83 45 C4 FC 03 46 C4 FB 93 07 B4 FA 03 47 D4 FE
83 46 E4 FE 13 05 C4 FA EF F0 5F DB 93 07 05 00
A3 0E F4 FC 03 47 D4 FD 93 07 10 00 63 14 F7 04
83 47 A4 FE 63 90 07 02 93 07 90 00 23 07 F4 FE
93 07 90 00 A3 06 F4 FE 93 07 10 00 23 05 F4 FE
6F 00 80 01 93 07 D0 01 23 07 F4 FE 93 07 D0 01
A3 06 F4 FE 23 05 04 FE 83 47 C4 FE 93 87 17 00
23 06 F4 FE 93 05 40 01 13 05 30 00 EF F0 8F 80
B7 07 40 00 13 85 C7 2D EF E0 5F DF 83 47 D4 FE
93 97 17 00 03 47 E4 FE 13 06 07 00 93 85 07 00
13 05 F0 04 EF E0 DF D0 93 06 C4 FB 13 06 C4 FC
93 05 C4 FA 83 47 D4 FD 13 07 F0 00 13 85 07 00
EF F0 5F BE 83 47 C4 FE 93 87 07 03 93 F7 F7 0F
13 06 70 02 93 05 30 00 13 85 07 00 EF E0 5F CD
83 47 C4 FC 63 82 07 02 03 47 C4 FC 93 07 F0 04
63 0C F7 00 83 47 C4 FB 63 88 07 00 03 47 C4 FB
93 07 B0 03 63 16 F7 00 93 07 10 00 6F 00 80 00
93 07 00 00 A3 05 F4 FE A3 0E 04 FC EF F0 0F 81
6F F0 1F D7 13 01 01 F7 23 26 11 08 23 24 81 08
13 04 01 09 EF E0 5F F9 B7 07 C0 00 83 A7 07 00
23 24 F4 FC 93 07 20 01 23 22 F4 FC 83 27 84 FC
93 87 C7 FF 13 07 70 00 E3 6C F7 1E 13 97 27 00
B7 07 40 00 93 87 C7 50 B3 07 F7 00 83 A7 07 00
67 80 07 00 B7 07 C0 01 93 87 07 15 23 A0 07 00
EF E0 DF FA 93 05 10 00 13 05 E0 01 EF E0 9F EF
B7 07 40 00 13 85 87 2E EF E0 5F CE B7 07 40 00
13 87 C7 3E 93 07 84 F7 93 06 07 00 13 07 80 04
13 06 07 00 93 85 06 00 13 85 07 00 EF 00 50 1B
23 24 04 FE 6F 00 C0 03 83 27 84 FE 93 97 27 00
13 07 04 FF B3 07 F7 00 03 A7 87 F8 B7 17 00 00
93 86 07 E1 13 06 00 00 83 25 84 FE 13 05 07 00
EF E0 1F F8 83 27 84 FE 93 87 17 00 23 24 F4 FE
03 27 84 FE 83 27 44 FC E3 40 F7 FC EF E0 1F F2
13 07 84 F7 B7 17 00 00 93 86 07 E1 13 06 00 00
83 25 44 FC 13 05 07 00 EF F0 4F 88 EF E0 1F F0
6F 00 00 00 EF F0 CF B2 23 20 04 FC B7 27 C0 03
93 87 47 02 83 A7 07 00 23 20 F4 FC 03 27 04 FC
93 07 10 00 63 14 F7 04 13 06 20 01 93 05 80 02
13 05 10 00 EF E0 9F D5 13 06 20 01 93 05 20 03
13 05 50 00 EF E0 9F D4 13 06 20 01 93 05 C0 03
13 05 50 00 EF E0 9F D3 13 06 20 01 93 05 60 04
13 05 50 00 EF E0 9F D2 6F F0 5F FA 03 27 04 FC
93 07 20 00 63 14 F7 04 13 06 20 01 93 05 20 03
13 05 10 00 EF E0 9F D0 13 06 20 01 93 05 80 02
13 05 50 00 EF E0 9F CF 13 06 20 01 93 05 C0 03
13 05 50 00 EF E0 9F CE 13 06 20 01 93 05 60 04
13 05 50 00 EF E0 9F CD 6F F0 5F F5 03 27 04 FC
93 07 40 00 63 14 F7 04 13 06 20 01 93 05 C0 03
13 05 10 00 EF E0 9F CB 13 06 20 01 93 05 80 02
13 05 50 00 EF E0 9F CA 13 06 20 01 93 05 20 03
13 05 50 00 EF E0 9F C9 13 06 20 01 93 05 60 04
13 05 50 00 EF E0 9F C8 6F F0 5F F0 03 27 04 FC
93 07 50 00 63 14 F7 04 13 06 20 01 93 05 60 04
13 05 10 00 EF E0 9F C6 13 06 20 01 93 05 80 02
13 05 50 00 EF E0 9F C5 13 06 20 01 93 05 20 03
13 05 50 00 EF E0 9F C4 13 06 20 01 93 05 C0 03
13 05 50 00 EF E0 9F C3 6F F0 5F EB 03 27 04 FC
93 07 10 08 63 06 F7 06 03 27 04 FC 93 07 20 08
63 00 F7 06 03 27 04 FC 93 07 40 08 63 0A F7 04
03 27 04 FC 93 07 50 08 63 04 F7 04 13 06 20 01
93 05 80 02 13 05 50 00 EF E0 5F BF 13 06 20 01
93 05 20 03 13 05 50 00 EF E0 5F BE 13 06 20 01
93 05 C0 03 13 05 50 00 EF E0 5F BD 13 06 20 01
93 05 60 04 13 05 50 00 EF E0 5F BC 6F F0 1F E4
03 27 04 FC 93 07 10 08 63 18 F7 00 EF E0 DF CB
EF F0 8F C7 6F 00 00 00 03 27 04 FC 93 07 20 08
63 18 F7 00 EF E0 5F CA EF F0 4F A0 6F 00 00 00
03 27 04 FC 93 07 50 08 63 18 F7 00 EF E0 DF C8
EF F0 DF A1 6F 00 00 00 03 27 04 FC 93 07 40 08
63 12 F7 70 EF E0 5F C7 B7 07 C0 02 13 87 C7 15
93 07 10 00 23 20 F7 00 37 07 C0 02 13 07 87 15
23 20 F7 00 37 07 C0 02 13 07 47 15 23 20 F7 00
37 07 C0 02 13 07 07 15 23 20 F7 00 37 07 C0 01
13 07 C7 15 23 20 F7 00 37 07 C0 01 13 07 87 15
23 20 F7 00 37 07 C0 01 13 07 07 15 23 20 F7 00
EF E0 DF C7 93 05 80 02 13 05 A0 05 EF E0 9F BC
B7 07 40 00 13 85 47 30 EF E0 5F 9B B7 07 40 00
13 87 47 43 93 07 84 F7 93 06 07 00 13 07 80 04
13 06 07 00 93 85 06 00 13 85 07 00 EF 00 40 68
23 22 04 FE 6F 00 00 04 83 27 44 FE 93 97 27 00
13 07 04 FF B3 07 F7 00 03 A7 87 F8 B7 17 00 00
93 86 07 E1 B7 17 00 00 13 86 87 2E 83 25 44 FE
13 05 07 00 EF E0 DF C4 83 27 44 FE 93 87 17 00
23 22 F4 FE 03 27 44 FE 83 27 44 FC E3 4E F7 FA
EF E0 DF BE 13 07 84 F7 B7 17 00 00 93 86 07 E1
B7 17 00 00 13 86 87 2E 83 25 44 FC 13 05 07 00
EF E0 DF D4 EF E0 9F BC 6F 00 00 00 B7 07 C0 01
93 87 87 15 23 A0 07 00 23 26 04 FE 6F 00 C0 0B
83 27 C4 FE 13 97 27 00 B7 07 40 03 B3 07 F7 00
13 07 F0 FF 23 A0 E7 00 03 27 C4 FE B7 17 00 00
93 87 07 96 B3 07 F7 00 13 97 27 00 B7 07 40 03
93 87 07 EC B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
03 27 C4 FE B7 17 00 00 93 87 07 2C B3 07 F7 00
13 97 27 00 B7 07 40 03 93 87 07 EC B3 07 F7 00
13 07 F0 FF 23 A0 E7 00 03 27 C4 FE B7 27 00 00
93 87 07 C2 B3 07 F7 00 13 97 27 00 B7 07 40 03
93 87 07 EC B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
83 27 C4 FE 13 97 27 00 B7 97 40 03 93 87 07 4C
B3 07 F7 00 13 07 F0 FF 23 A0 E7 00 83 27 C4 FE
93 87 17 00 23 26 F4 FE 03 27 C4 FE 93 07 F0 04
E3 D0 E7 F4 23 26 04 FE 6F 00 00 09 03 27 C4 FE
93 07 07 00 93 97 27 00 B3 87 E7 00 93 97 67 00
13 87 07 00 B7 07 40 03 B3 07 F7 00 13 07 F0 FF
23 A0 E7 00 03 27 C4 FE 93 07 07 00 93 97 27 00
B3 87 E7 00 93 97 67 00 13 87 07 00 B7 07 40 03
93 87 C7 09 B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
03 27 C4 FE 93 07 07 00 93 97 27 00 B3 87 E7 00
93 97 67 00 13 87 07 00 B7 07 40 03 93 87 C7 13
B3 07 F7 00 13 07 F0 FF 23 A0 E7 00 83 27 C4 FE
93 87 17 00 23 26 F4 FE 03 27 C4 FE 93 07 70 07
E3 D6 E7 F6 EF E0 9F A4 93 05 80 02 13 05 E0 01
EF E0 5F 99 B7 07 40 00 13 85 47 32 EF E0 0F F8
B7 07 40 00 13 87 C7 47 93 07 84 F7 93 06 07 00
13 07 80 04 13 06 07 00 93 85 06 00 13 85 07 00
EF 00 00 45 23 20 04 FE 6F 00 C0 03 83 27 04 FE
93 97 27 00 13 07 04 FF B3 07 F7 00 03 A7 87 F8
B7 17 00 00 93 86 07 E1 13 06 80 02 83 25 04 FE
13 05 07 00 EF E0 DF A1 83 27 04 FE 93 87 17 00
23 20 F4 FE 03 27 04 FE 83 27 44 FC E3 40 F7 FC
EF E0 DF 9B 13 07 84 F7 B7 17 00 00 93 86 07 E1
13 06 80 02 83 25 44 FC 13 05 07 00 EF E0 1F B2
EF E0 DF 99 6F 00 00 00 B7 07 C0 01 93 87 C7 15
23 A0 07 00 EF E0 9F 98 93 05 10 00 13 05 A0 05
EF E0 5F 8D B7 07 40 00 13 85 07 34 EF E0 0F EC
B7 07 40 00 13 87 47 4C 93 07 84 F7 93 06 07 00
13 07 80 04 13 06 07 00 93 85 06 00 13 85 07 00
EF 00 00 39 23 2E 04 FC 6F 00 00 04 83 27 C4 FD
93 97 27 00 13 07 04 FF B3 07 F7 00 03 A7 87 F8
B7 17 00 00 93 86 07 E1 B7 17 00 00 13 86 07 2C
83 25 C4 FD 13 05 07 00 EF E0 9F 95 83 27 C4 FD
93 87 17 00 23 2E F4 FC 03 27 C4 FD 83 27 44 FC
E3 4E F7 FA EF E0 9F 8F 13 07 84 F7 B7 17 00 00
93 86 07 E1 B7 17 00 00 13 86 07 2C 83 25 44 FC
13 05 07 00 EF E0 9F A5 EF E0 5F 8D 6F 00 00 00
B7 07 C0 02 93 87 07 15 23 A0 07 00 EF E0 1F 8C
93 05 10 00 13 05 10 00 EF E0 DF 80 B7 07 40 00
13 85 47 36 EF E0 8F DF B7 07 40 00 13 87 C7 3E
93 07 84 F7 93 06 07 00 13 07 80 04 13 06 07 00
93 85 06 00 13 85 07 00 EF 00 80 2C 23 2C 04 FC
6F 00 80 03 83 27 84 FD 93 97 27 00 13 07 04 FF
B3 07 F7 00 83 A7 87 F8 93 06 00 4B 13 06 00 00
83 25 84 FD 13 85 07 00 EF E0 9F 89 83 27 84 FD
93 87 17 00 23 2C F4 FC 03 27 84 FD 83 27 44 FC
E3 42 F7 FC EF E0 9F 83 93 07 84 F7 93 06 00 4B
13 06 00 00 83 25 44 FC 13 85 07 00 EF E0 9F AE
EF E0 DF 81 6F 00 00 00 B7 07 C0 02 93 87 47 15
23 A0 07 00 EF E0 9F 80 93 05 80 02 13 05 C0 03
EF E0 4F F5 B7 07 40 00 13 85 47 38 EF E0 0F D4
B7 07 40 00 13 87 47 43 93 07 84 F7 93 06 07 00
13 07 80 04 13 06 07 00 93 85 06 00 13 85 07 00
EF 00 00 21 23 2A 04 FC 6F 00 C0 03 83 27 44 FD
93 97 27 00 13 07 04 FF B3 07 F7 00 03 A7 87 F8
93 06 00 4B B7 17 00 00 13 86 87 2E 83 25 44 FD
13 05 07 00 EF E0 CF FD 83 27 44 FD 93 87 17 00
23 2A F4 FC 03 27 44 FD 83 27 44 FC E3 40 F7 FC
EF E0 CF F7 13 07 84 F7 93 06 00 4B B7 17 00 00
13 86 87 2E 83 25 44 FC 13 05 07 00 EF E0 9F A2
EF E0 CF F5 6F 00 00 00 B7 07 C0 02 93 87 87 15
23 A0 07 00 EF E0 8F F4 93 05 80 02 13 05 10 00
EF E0 4F E9 B7 07 40 00 13 85 47 3A EF E0 0F C8
B7 07 40 00 13 87 C7 47 93 07 84 F7 93 06 07 00
13 07 80 04 13 06 07 00 93 85 06 00 13 85 07 00
EF 00 00 15 23 28 04 FC 6F 00 80 03 83 27 04 FD
93 97 27 00 13 07 04 FF B3 07 F7 00 83 A7 87 F8
93 06 00 4B 13 06 80 02 83 25 04 FD 13 85 07 00
EF E0 0F F2 83 27 04 FD 93 87 17 00 23 28 F4 FC
03 27 04 FD 83 27 44 FC E3 42 F7 FC EF E0 0F EC
93 07 84 F7 93 06 00 4B 13 06 80 02 83 25 44 FC
13 85 07 00 EF E0 1F 97 EF E0 4F EA 6F 00 00 00
B7 07 C0 02 93 87 C7 15 23 A0 07 00 EF E0 0F E9
93 05 10 00 13 05 C0 03 EF E0 CF DD B7 07 40 00
13 85 47 3C EF E0 8F BC B7 07 40 00 13 87 47 4C
93 07 84 F7 93 06 07 00 13 07 80 04 13 06 07 00
93 85 06 00 13 85 07 00 EF 00 80 09 23 26 04 FC
6F 00 C0 03 83 27 C4 FC 93 97 27 00 13 07 04 FF
B3 07 F7 00 03 A7 87 F8 93 06 00 4B B7 17 00 00
13 86 07 2C 83 25 C4 FC 13 05 07 00 EF E0 4F E6
83 27 C4 FC 93 87 17 00 23 26 F4 FC 03 27 C4 FC
83 27 44 FC E3 40 F7 FC EF E0 4F E0 13 07 84 F7
93 06 00 4B B7 17 00 00 13 86 07 2C 83 25 44 FC
13 05 07 00 EF E0 1F 8B EF E0 4F DE 6F 00 00 00
6F 00 00 00 13 00 00 00 93 07 00 00 13 85 07 00
83 20 C1 08 03 24 81 08 13 01 01 09 67 80 00 00
@00001E68
B3 C7 A5 00 93 F7 37 00 B3 08 C5 00 63 96 07 06
93 07 30 00 63 F2 C7 06 93 77 35 00 13 07 05 00
63 9A 07 0C 13 F6 C8 FF B3 06 E6 40 93 07 00 02
93 02 00 02 63 C2 D7 06 93 86 05 00 93 07 07 00
63 78 C7 02 03 A8 06 00 93 87 47 00 93 86 46 00
23 AE 07 FF E3 E8 C7 FE 93 07 F6 FF B3 87 E7 40
93 F7 C7 FF 93 87 47 00 33 07 F7 00 B3 85 F5 00
63 68 17 01 67 80 00 00 13 07 05 00 E3 7C 15 FF
83 C7 05 00 13 07 17 00 93 85 15 00 A3 0F F7 FE
E3 68 17 FF 67 80 00 00 83 A6 45 00 83 A7 C5 01
83 AF 05 00 03 AF 85 00 83 AE C5 00 03 AE 05 01
03 A3 45 01 03 A8 85 01 23 22 D7 00 83 A6 05 02
23 20 F7 01 23 24 E7 01 23 26 D7 01 23 28 C7 01
23 2A 67 00 23 2C 07 01 23 2E F7 00 13 07 47 02
B3 07 E6 40 23 2E D7 FE 93 85 45 02 E3 C6 F2 FA
6F F0 9F F4 83 C6 05 00 13 07 17 00 93 77 37 00
A3 0F D7 FE 93 85 15 00 E3 8E 07 F0 83 C6 05 00
13 07 17 00 93 77 37 00 A3 0F D7 FE 93 85 15 00
E3 9A 07 FC 6F F0 1F F0
