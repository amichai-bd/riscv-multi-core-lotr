/*
 RC to wishbone gateway controller
 this module controlls the uart ip 
 via wishbone transactions and the 
 lotr project via the RC controller
 */

`timescale 1ns/1ns

module gateway
  #()
   (
    // RC Interface
    // wishbone interface
    );

endmodule // gateway
