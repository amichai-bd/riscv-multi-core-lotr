@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 93 00 00 00 13 01 00 00 93 01 00 00
13 02 00 00 93 02 00 00 13 03 00 00 93 03 00 00
13 04 00 00 93 04 00 00 13 05 00 00 93 05 00 00
13 06 00 00 93 06 00 00 13 07 00 00 93 07 00 00
13 08 00 00 93 08 00 00 13 09 00 00 93 09 00 00
13 0A 00 00 93 0A 00 00 13 0B 00 00 93 0B 00 00
13 0C 00 00 93 0C 00 00 13 0D 00 00 93 0D 00 00
13 0E 00 00 93 0E 00 00 13 0F 00 00 93 0F 00 00
B7 02 C0 00 83 A2 42 00 93 05 00 07 13 86 12 00
EF 00 80 0C 37 06 40 00 13 06 06 64 33 01 C5 00
13 04 01 00 93 05 00 02 13 86 02 00 EF 00 C0 0A
B7 06 40 00 B3 86 A6 00 23 A0 56 00 37 03 40 00
13 03 03 08 23 A2 66 00 13 03 00 08 23 A4 66 00
93 05 00 15 13 86 02 00 EF 00 00 08 37 03 40 00
13 03 03 10 33 03 A3 00 23 A6 66 00 13 03 00 15
23 A8 66 00 13 03 40 01 93 03 00 02 33 85 66 00
23 20 05 00 13 03 43 00 E3 4A 73 FE 83 A1 46 00
03 A2 C6 00 93 03 00 00 63 8A 72 00 37 03 C0 00
83 23 03 20 E3 8C 03 FE 6F 00 80 01 13 85 06 00
EF 00 00 04 37 03 C0 00 93 03 10 00 23 20 73 20
13 85 06 00 EF 00 40 06 13 85 06 00 EF 00 80 0C
6F F0 9F FF 73 00 10 00 13 05 00 00 63 08 06 00
33 05 B5 00 13 06 F6 FF E3 1C 06 FE 67 80 00 00
13 01 01 FF 23 24 81 00 03 24 45 00 13 06 00 00
93 05 40 01 13 05 04 00 23 26 11 00 EF 00 00 16
93 07 50 3E 83 20 C1 00 23 20 F4 00 03 24 81 00
13 01 01 01 67 80 00 00 13 01 01 FF 23 22 91 00
83 24 C5 00 23 24 81 00 13 06 00 00 13 04 05 00
93 05 80 00 13 85 04 00 23 20 21 01 23 26 11 00
03 29 44 00 EF 00 80 11 03 27 04 00 63 00 07 02
83 27 09 00 93 06 30 00 23 A2 D4 00 93 D7 17 00
B3 87 E7 40 93 87 17 00 23 A0 F4 00 83 20 C1 00
03 24 81 00 83 24 41 00 03 29 01 00 13 01 01 01
67 80 00 00 83 27 05 00 03 26 45 00 63 9E 07 04
83 27 C6 00 83 26 86 00 03 27 06 01 93 F5 17 00
93 F6 36 00 B3 E6 B6 00 93 F7 27 00 93 75 17 00
93 C6 16 00 B3 E6 D7 00 93 C7 F5 FF B3 F6 D7 00
83 25 46 00 93 77 27 00 B3 E7 D7 00 13 F7 27 00
93 C7 F7 FF 33 67 B7 00 93 F7 17 00 B3 67 F7 00
23 22 F6 00 67 80 00 00 03 25 C5 00 93 97 27 00
B3 06 F6 00 03 27 05 00 93 07 10 00 83 A5 46 00
63 FA E7 02 93 F7 15 00 63 98 07 04 83 27 06 00
63 78 F7 02 B3 87 E7 40 E3 6E F7 FE 83 27 45 00
93 E5 35 00 23 A2 B6 00 63 72 F7 02 23 20 05 00
67 80 00 00 93 E5 15 00 23 A2 B6 00 67 80 00 00
E3 9E 07 FC 83 27 45 00 E3 62 F7 FE 33 07 F7 40
23 20 E5 00 67 80 00 00 67 80 00 00 63 8A 05 00
B3 05 B5 00 23 20 C5 00 13 05 45 00 E3 1C B5 FE
67 80 00 00 83 27 05 00 E3 8E 07 FE 03 25 05 00
67 80 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
