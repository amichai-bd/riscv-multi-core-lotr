@00400000
0B 00 00 00 05 00 00 00 09 00 00 00 0D 00 00 00
12 00 00 00 07 00 00 00 01 00 00 00 02 00 00 00
0C 00 00 00 0A 00 00 00 04 00 00 00 03 00 00 00
0E 00 00 00 06 00 00 00 0F 00 00 00 11 00 00 00
08 00 00 00 10 00 00 00 01 00 00 00 02 00 00 00
03 00 00 00 04 00 00 00 05 00 00 00 06 00 00 00
0D 00 00 00 0E 00 00 00 0F 00 00 00 10 00 00 00
11 00 00 00 12 00 00 00 07 00 00 00 08 00 00 00
09 00 00 00 0A 00 00 00 0B 00 00 00 0C 00 00 00
12 00 00 00 11 00 00 00 10 00 00 00 0F 00 00 00
0E 00 00 00 0D 00 00 00 0C 00 00 00 0B 00 00 00
0A 00 00 00 09 00 00 00 08 00 00 00 07 00 00 00
06 00 00 00 05 00 00 00 04 00 00 00 03 00 00 00
02 00 00 00 01 00 00 00 02 00 00 00 03 00 00 00
04 00 00 00 05 00 00 00 06 00 00 00 07 00 00 00
08 00 00 00 09 00 00 00 0A 00 00 00 0B 00 00 00
0C 00 00 00 0D 00 00 00 0E 00 00 00 0F 00 00 00
10 00 00 00 11 00 00 00 12 00 00 00 01 00 00 00
20 05 00 00 C4 05 00 00 70 06 00 00 80 08 00 00
2C 09 00 00 C8 09 00 00 6C 0A 00 00 08 0B 00 00
