@00400800
3C 0C 00 00 50 0C 00 00 5C 0C 00 00 68 0C 00 00
74 0C 00 00 80 0C 00 00 8C 0C 00 00 98 0C 00 00
