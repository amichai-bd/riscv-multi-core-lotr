@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
6F 00 00 32 67 80 00 00
@00000088
13 01 01 FD 23 26 11 02 23 24 81 02 23 22 91 02
13 04 01 03 23 2E A4 FC 23 2C B4 FC 23 2A C4 FC
23 26 04 FE 6F 00 80 15 23 24 04 FE 6F 00 80 13
03 27 C4 FE 93 07 07 00 93 97 17 00 B3 87 E7 00
93 97 27 00 13 87 07 00 83 27 44 FD 33 87 E7 00
83 27 84 FE 93 97 27 00 B3 07 F7 00 23 A0 07 00
23 22 04 FE 6F 00 80 0E 03 27 C4 FE 93 07 07 00
93 97 17 00 B3 87 E7 00 93 97 27 00 13 87 07 00
83 27 44 FD 33 87 E7 00 83 27 84 FE 93 97 27 00
B3 07 F7 00 83 A4 07 00 03 27 C4 FE 93 07 07 00
93 97 17 00 B3 87 E7 00 93 97 27 00 13 87 07 00
83 27 C4 FD 33 87 E7 00 83 27 44 FE 93 97 27 00
B3 07 F7 00 83 A6 07 00 03 27 44 FE 93 07 07 00
93 97 17 00 B3 87 E7 00 93 97 27 00 13 87 07 00
83 27 84 FD 33 87 E7 00 83 27 84 FE 93 97 27 00
B3 07 F7 00 83 A7 07 00 93 85 07 00 13 85 06 00
EF 00 80 26 93 07 05 00 13 86 07 00 03 27 C4 FE
93 07 07 00 93 97 17 00 B3 87 E7 00 93 97 27 00
13 87 07 00 83 27 44 FD B3 86 E7 00 33 87 C4 00
83 27 84 FE 93 97 27 00 B3 87 F6 00 23 A0 E7 00
83 27 44 FE 93 87 17 00 23 22 F4 FE 03 27 44 FE
93 07 20 00 E3 DA E7 F0 83 27 84 FE 93 87 17 00
23 24 F4 FE 03 27 84 FE 93 07 20 00 E3 D2 E7 EC
83 27 C4 FE 93 87 17 00 23 26 F4 FE 03 27 C4 FE
93 07 20 00 E3 D2 E7 EA 13 00 00 00 13 00 00 00
83 20 C1 02 03 24 81 02 83 24 41 02 13 01 01 03
67 80 00 00 13 01 01 F8 23 2E 11 06 23 2C 81 06
13 04 01 08 93 07 10 00 23 26 F4 FC 93 07 20 00
23 28 F4 FC 93 07 30 00 23 2A F4 FC 93 07 40 00
23 2C F4 FC 93 07 50 00 23 2E F4 FC 93 07 60 00
23 20 F4 FE 93 07 70 00 23 22 F4 FE 93 07 80 00
23 24 F4 FE 93 07 90 00 23 26 F4 FE 93 07 90 00
23 24 F4 FA 93 07 80 00 23 26 F4 FA 93 07 70 00
23 28 F4 FA 93 07 60 00 23 2A F4 FA 93 07 50 00
23 2C F4 FA 93 07 40 00 23 2E F4 FA 93 07 30 00
23 20 F4 FC 93 07 20 00 23 22 F4 FC 93 07 10 00
23 24 F4 FC 93 06 44 F8 13 07 84 FA 93 07 C4 FC
13 86 06 00 93 05 07 00 13 85 07 00 EF F0 5F DA
B7 17 40 00 93 87 07 F0 03 27 44 F8 23 A0 E7 00
B7 17 40 00 93 87 07 F0 03 27 84 F8 23 A2 E7 00
B7 17 40 00 93 87 07 F0 03 27 C4 F8 23 A4 E7 00
B7 17 40 00 93 87 07 F0 03 27 04 F9 23 A6 E7 00
B7 17 40 00 93 87 07 F0 03 27 44 F9 23 A8 E7 00
B7 17 40 00 93 87 07 F0 03 27 84 F9 23 AA E7 00
B7 17 40 00 93 87 07 F0 03 27 C4 F9 23 AC E7 00
B7 17 40 00 93 87 07 F0 03 27 04 FA 23 AE E7 00
B7 17 40 00 93 87 07 F0 03 27 44 FA 23 A0 E7 02
B7 17 40 00 93 87 07 F0 13 07 F0 0F 23 AE E7 0E
93 07 00 00 13 85 07 00 83 20 C1 07 03 24 81 07
13 01 01 08 67 80 00 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 17 11 40 00 13 01 41 B2 13 05 00 00
93 05 00 00 EF F0 1F E4 13 06 05 00 13 05 00 00
93 F6 15 00 63 84 06 00 33 05 C5 00 93 D5 15 00
13 16 16 00 E3 96 05 FE 67 80 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00
