@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 80 00 73 00 10 00
@000000A8
13 01 01 B2 23 2E 11 4C 23 2C 81 4C 13 04 01 4E
B7 07 C0 00 93 87 47 00 83 A7 07 00 23 22 F4 FE
B7 07 C0 00 93 87 87 00 83 A7 07 00 23 20 F4 FE
B7 07 40 00 13 87 07 00 93 07 84 D9 93 06 07 00
13 07 00 24 13 06 07 00 93 85 06 00 13 85 07 00
EF 00 80 27 B7 07 40 00 13 87 07 24 93 07 84 B5
93 06 07 00 13 07 00 24 13 06 07 00 93 85 06 00
13 85 07 00 EF 00 40 25 83 27 04 FE 13 97 27 00
83 27 44 FE 33 07 F7 00 93 06 84 D9 93 07 07 00
93 97 17 00 B3 87 E7 00 93 97 47 00 B3 87 F6 00
23 2E F4 FC 83 27 04 FE 13 97 27 00 83 27 44 FE
33 07 F7 00 93 06 84 B5 93 07 07 00 93 97 17 00
B3 87 E7 00 93 97 47 00 B3 87 F6 00 23 2C F4 FC
23 26 04 FE 6F 00 00 06 83 27 C4 FE 93 97 27 00
03 27 C4 FD B3 07 F7 00 83 A6 07 00 83 27 C4 FE
93 97 27 00 03 27 84 FD B3 07 F7 00 83 A7 07 00
93 85 07 00 13 85 06 00 EF 00 C0 19 93 07 05 00
13 87 07 00 83 27 C4 FE 93 97 27 00 93 87 07 FF
B3 87 87 00 23 AC E7 B2 83 27 C4 FE 93 87 17 00
23 26 F4 FE 03 27 C4 FE 93 07 B0 00 E3 DE E7 F8
23 24 04 FE 6F 00 40 06 83 27 04 FE 13 97 27 00
83 27 44 FE 33 07 F7 00 93 07 07 00 93 97 17 00
B3 87 E7 00 93 97 27 00 13 87 07 00 83 27 84 FE
B3 07 F7 00 13 97 27 00 B7 17 40 01 93 87 07 F0
33 07 F7 00 83 27 84 FE 93 97 27 00 93 87 07 FF
B3 87 87 00 83 A7 87 B3 23 20 F7 00 83 27 84 FE
93 87 17 00 23 24 F4 FE 03 27 84 FE 93 07 B0 00
E3 DC E7 F8 83 27 44 FE 63 84 07 02 03 27 04 FE
93 07 10 00 63 0E F7 00 83 27 44 FE 93 97 27 00
93 87 07 20 13 07 10 00 23 A0 E7 00 6F 00 00 00
03 27 04 FE 93 07 10 00 63 06 F7 04 13 00 00 00
93 07 40 20 83 A7 07 00 E3 8C 07 FE 93 07 80 20
83 A7 07 00 E3 86 07 FE 93 07 C0 20 83 A7 07 00
E3 80 07 FE 83 27 04 FE 13 97 27 00 B7 07 00 01
93 87 07 20 B3 07 F7 00 13 07 10 00 23 A0 E7 00
6F 00 C0 05 83 27 44 FE 63 8E 07 00 93 07 40 20
03 A7 07 00 93 07 40 20 13 07 17 00 23 A0 E7 00
6F 00 00 00 13 00 00 00 93 07 00 20 83 A7 07 00
E3 8C 07 FE 93 07 80 20 83 A7 07 00 E3 86 07 FE
93 07 C0 20 83 A7 07 00 E3 80 07 FE 93 07 40 20
03 A7 07 00 93 07 30 00 E3 18 F7 FC 13 00 00 00
13 85 07 00 83 20 C1 4D 03 24 81 4D 13 01 01 4E
67 80 00 00 13 06 05 00 13 05 00 00 93 F6 15 00
63 84 06 00 33 05 C5 00 93 D5 15 00 13 16 16 00
E3 96 05 FE 67 80 00 00 B3 47 B5 00 93 F7 37 00
B3 08 C5 00 63 96 07 06 93 07 30 00 63 F2 C7 06
93 77 35 00 13 07 05 00 63 9A 07 0C 13 F6 C8 FF
B3 06 E6 40 93 07 00 02 93 02 00 02 63 C2 D7 06
93 86 05 00 93 07 07 00 63 78 C7 02 03 A8 06 00
93 87 47 00 93 86 46 00 23 AE 07 FF E3 E8 C7 FE
93 07 F6 FF B3 87 E7 40 93 F7 C7 FF 93 87 47 00
33 07 F7 00 B3 85 F5 00 63 68 17 01 67 80 00 00
13 07 05 00 E3 7C 15 FF 83 C7 05 00 13 07 17 00
93 85 15 00 A3 0F F7 FE E3 68 17 FF 67 80 00 00
83 A6 45 00 83 A7 C5 01 83 AF 05 00 03 AF 85 00
83 AE C5 00 03 AE 05 01 03 A3 45 01 03 A8 85 01
23 22 D7 00 83 A6 05 02 23 20 F7 01 23 24 E7 01
23 26 D7 01 23 28 C7 01 23 2A 67 00 23 2C 07 01
23 2E F7 00 13 07 47 02 B3 07 E6 40 23 2E D7 FE
93 85 45 02 E3 C6 F2 FA 6F F0 9F F4 83 C6 05 00
13 07 17 00 93 77 37 00 A3 0F D7 FE 93 85 15 00
E3 8E 07 F0 83 C6 05 00 13 07 17 00 93 77 37 00
A3 0F D7 FE 93 85 15 00 E3 9A 07 FC 6F F0 1F F0
