@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 80 00 73 00 10 00
@000000A8
13 01 01 FE 23 2E 11 00 23 2C 81 00 23 2A 91 00
13 04 01 02 B7 07 C0 00 83 A7 07 00 23 26 F4 FE
03 27 C4 FE 93 07 40 00 63 1A F7 06 B7 17 40 00
83 A7 07 80 23 24 F4 FE B7 17 40 00 83 A7 47 80
23 22 F4 FE B7 17 40 00 93 84 07 F0 83 25 44 FE
03 25 84 FE EF 00 80 06 93 07 05 00 23 A0 F4 00
B7 17 40 00 93 84 47 F0 83 25 44 FE 03 25 84 FE
EF 00 D0 03 93 07 05 00 23 A0 F4 00 B7 17 40 00
93 84 87 F0 83 25 84 FE 03 25 44 FE EF 00 C0 48
93 07 05 00 23 A0 F4 00 6F 00 80 00 6F 00 00 00
93 07 00 00 13 85 07 00 83 20 C1 01 03 24 81 01
83 24 41 01 13 01 01 02 67 80 00 00 37 07 80 00
13 01 01 FF 13 07 F7 FF B3 77 A7 00 23 24 81 00
23 22 91 00 13 54 75 01 93 54 F5 01 13 D5 75 01
33 77 B7 00 13 74 F4 0F 13 75 F5 0F 23 26 11 00
23 20 21 01 93 D5 F5 01 93 97 37 00 13 17 37 00
B3 06 A4 40 63 9A B4 18 63 50 D0 0A 63 16 05 02
63 00 07 18 13 86 F6 FF 63 18 06 00 B3 87 E7 00
13 04 10 00 6F 00 00 05 93 05 F0 0F 63 90 B6 02
13 04 F0 0F 6F 00 80 11 13 06 F0 0F 63 08 C4 10
37 06 00 04 33 67 C7 00 13 86 06 00 93 05 B0 01
93 06 10 00 63 CE C5 00 93 06 00 02 B3 86 C6 40
B3 55 C7 00 33 17 D7 00 33 37 E0 00 B3 E6 E5 00
B3 87 D7 00 37 07 00 04 33 F7 E7 00 63 08 07 0C
13 04 14 00 13 07 F0 0F 63 02 E4 30 37 07 00 7E
93 F6 17 00 13 07 F7 FF 93 D7 17 00 B3 F7 E7 00
B3 E7 D7 00 6F 00 80 0A 63 86 06 06 B3 06 85 40
63 10 04 02 63 82 07 2C 13 86 F6 FF E3 00 06 F6
93 05 F0 0F 63 90 B6 02 93 07 07 00 6F F0 5F F6
13 06 F0 0F E3 0A C5 FE 37 06 00 04 B3 E7 C7 00
13 86 06 00 93 05 B0 01 93 06 10 00 63 CE C5 00
93 06 00 02 B3 86 C6 40 B3 D5 C7 00 B3 97 D7 00
B3 37 F0 00 B3 E6 F5 00 B3 87 E6 00 13 04 05 00
6F F0 5F F6 93 06 14 00 13 F6 E6 0F 63 12 06 06
63 14 04 04 63 8E 07 24 63 02 07 02 B3 87 E7 00
37 07 00 04 33 F7 E7 00 63 0A 07 00 37 07 00 FC
13 07 F7 FF B3 F7 E7 00 13 04 10 00 13 F7 77 00
63 00 07 24 13 F7 F7 00 93 06 40 00 63 0A D7 22
93 87 47 00 6F 00 C0 22 E3 80 07 F6 E3 02 07 EC
93 04 00 00 B7 07 00 02 13 04 F0 0F 6F 00 40 21
13 06 F0 0F 63 82 C6 20 B3 87 E7 00 93 D7 17 00
13 84 06 00 6F F0 9F FB 63 50 D0 08 63 12 05 06
E3 08 07 FE 13 86 F6 FF 63 18 06 00 B3 87 E7 40
13 04 10 00 6F 00 40 03 93 05 F0 0F E3 8A B6 E6
93 05 B0 01 93 06 10 00 63 CE C5 00 93 06 00 02
B3 86 C6 40 B3 55 C7 00 33 17 D7 00 33 37 E0 00
B3 E6 E5 00 B3 87 D7 40 37 09 00 04 33 F7 27 01
E3 0E 07 F4 13 09 F9 FF 33 F9 27 01 6F 00 80 11
13 06 F0 0F E3 04 C4 F4 37 06 00 04 33 67 C7 00
13 86 06 00 6F F0 DF FA 63 80 06 08 B3 06 85 40
63 18 04 02 63 80 07 1E 13 86 F6 FF 63 18 06 00
B3 07 F7 40 93 84 05 00 6F F0 9F F7 13 08 F0 0F
63 92 06 03 93 07 07 00 13 04 F0 0F 6F 00 C0 06
13 06 F0 0F E3 08 C5 FE 37 06 00 04 B3 E7 C7 00
13 86 06 00 13 08 B0 01 93 06 10 00 63 4E C8 00
93 06 00 02 B3 86 C6 40 33 D8 C7 00 B3 97 D7 00
B3 37 F0 00 B3 66 F8 00 B3 07 D7 40 13 04 05 00
93 84 05 00 6F F0 5F F5 93 06 14 00 93 F6 E6 0F
63 9E 06 04 63 12 04 04 63 9C 07 00 93 04 00 00
63 00 07 0E 93 07 07 00 93 84 05 00 6F F0 1F E9
E3 06 07 E8 B3 86 E7 40 37 06 00 04 33 F6 C6 00
B3 07 F7 40 E3 12 06 FE 93 07 00 00 63 80 06 08
93 87 06 00 6F F0 9F E6 E3 92 07 E8 E3 02 07 E8
93 07 07 00 93 84 05 00 6F F0 9F D3 33 89 E7 40
B7 06 00 04 B3 76 D9 00 63 84 06 04 33 09 F7 40
93 84 05 00 13 05 09 00 EF 00 D0 09 13 05 B5 FF
33 19 A9 00 63 40 85 04 33 05 85 40 13 05 15 00
13 04 00 02 B3 57 A9 00 33 05 A4 40 33 19 A9 00
33 39 20 01 B3 E7 27 01 13 04 00 00 6F F0 1F E0
E3 12 09 FC 93 07 00 00 13 04 00 00 93 04 00 00
6F 00 00 03 B7 07 00 FC 93 87 F7 FF 33 04 A4 40
B3 77 F9 00 6F F0 9F DD 93 07 07 00 6F F0 5F E1
93 07 07 00 6F F0 9F DC 13 04 F0 0F 93 07 00 00
37 07 00 04 33 F7 E7 00 63 0E 07 00 13 04 14 00
13 07 F0 0F 63 06 E4 06 37 07 00 FC 13 07 F7 FF
B3 F7 E7 00 13 07 F0 0F 93 D7 37 00 63 18 E4 00
63 86 07 00 B7 07 40 00 93 04 00 00 37 05 80 7F
13 14 74 01 93 97 97 00 33 74 A4 00 93 D7 97 00
83 20 C1 00 B3 67 F4 00 03 24 81 00 13 95 F4 01
03 29 01 00 83 24 41 00 33 E5 A7 00 13 01 01 01
67 80 00 00 93 07 07 00 13 84 06 00 6F F0 DF EA
93 07 00 00 6F F0 1F FA 13 01 01 FD 23 22 91 02
93 54 75 01 23 2E 31 01 23 2A 51 01 23 28 61 01
93 1A 95 00 23 26 11 02 23 24 81 02 23 20 21 03
23 2C 41 01 23 26 71 01 23 24 81 01 23 22 91 01
93 F4 F4 0F 13 8B 05 00 93 DA 9A 00 93 59 F5 01
63 84 04 08 93 07 F0 0F 63 80 F4 0A 93 9A 3A 00
B7 07 00 04 B3 EA FA 00 93 84 14 F8 93 0B 00 00
93 57 7B 01 13 14 9B 00 93 F7 F7 0F 13 54 94 00
13 5B FB 01 63 8A 07 08 13 07 F0 0F 63 86 E7 0A
13 14 34 00 37 07 00 04 33 64 E4 00 93 87 17 F8
13 07 00 00 93 96 2B 00 B3 E6 E6 00 33 8A F4 40
93 86 F6 FF 93 07 E0 00 33 C9 69 01 63 EE D7 08
B7 17 40 00 93 87 87 80 93 96 26 00 B3 86 F6 00
83 A7 06 00 67 80 07 00 63 8A 0A 02 13 85 0A 00
EF 00 40 6C 93 07 B5 FF 93 04 A0 F8 B3 9A FA 00
B3 84 A4 40 6F F0 9F F7 93 04 F0 0F 93 0B 20 00
E3 88 0A F6 93 0B 30 00 6F F0 9F F6 93 04 00 00
93 0B 10 00 6F F0 DF F5 63 0A 04 02 13 05 04 00
EF 00 40 68 93 07 B5 FF 33 14 F4 00 93 07 A0 F8
B3 87 A7 40 6F F0 DF F6 93 07 F0 0F 13 07 20 00
E3 02 04 F6 13 07 30 00 6F F0 DF F5 93 07 00 00
13 07 10 00 6F F0 1F F5 93 1C 54 00 63 FC 8A 16
13 0A FA FF 93 04 00 00 13 DB 0C 01 37 04 01 00
93 05 0B 00 13 04 F4 FF 13 85 0A 00 EF 00 C0 57
33 F4 8C 00 93 05 05 00 13 0C 05 00 13 05 04 00
EF 00 C0 53 93 0B 05 00 93 05 0B 00 13 85 0A 00
EF 00 00 5A 13 15 05 01 93 D7 04 01 B3 E7 A7 00
93 09 0C 00 63 FE 77 01 B3 87 97 01 93 09 FC FF
63 E8 97 01 63 F6 77 01 93 09 EC FF B3 87 97 01
B3 8B 77 41 93 05 0B 00 13 85 0B 00 EF 00 C0 51
93 05 05 00 93 0A 05 00 13 05 04 00 EF 00 00 4E
13 04 05 00 93 05 0B 00 13 85 0B 00 EF 00 40 54
93 17 05 01 13 87 0A 00 63 FE 87 00 B3 87 97 01
13 87 FA FF 63 E8 97 01 63 F6 87 00 13 87 EA FF
B3 87 97 01 B3 87 87 40 93 99 09 01 B3 E9 E9 00
B3 37 F0 00 33 E4 F9 00 13 07 FA 07 63 56 E0 0E
93 77 74 00 63 8A 07 00 93 77 F4 00 93 06 40 00
63 84 D7 00 13 04 44 00 B7 07 00 08 B3 77 F4 00
63 8A 07 00 B7 07 00 F8 93 87 F7 FF 33 74 F4 00
13 07 0A 08 93 07 E0 0F 13 54 34 00 63 C4 E7 08
93 17 77 01 13 14 94 00 37 07 80 7F B3 F7 E7 00
13 54 94 00 33 E4 87 00 13 15 F9 01 83 20 C1 02
33 65 A4 00 03 24 81 02 83 24 41 02 03 29 01 02
83 29 C1 01 03 2A 81 01 83 2A 41 01 03 2B 01 01
83 2B C1 00 03 2C 81 00 83 2C 41 00 13 01 01 03
67 80 00 00 93 94 FA 01 93 DA 1A 00 6F F0 DF E8
13 89 09 00 13 84 0A 00 13 87 0B 00 93 07 30 00
63 08 F7 08 93 07 10 00 63 0C F7 08 93 07 20 00
E3 1C F7 F2 13 04 00 00 13 07 F0 0F 6F F0 5F F7
13 09 0B 00 6F F0 9F FD 37 04 40 00 13 09 00 00
13 07 30 00 6F F0 9F FC 93 07 10 00 B3 87 E7 40
13 07 B0 01 63 4E F7 04 93 04 EA 09 B3 57 F4 00
33 14 94 00 33 34 80 00 33 E4 87 00 93 77 74 00
63 8A 07 00 93 77 F4 00 13 07 40 00 63 84 E7 00
13 04 44 00 B7 07 00 04 B3 77 F4 00 13 54 34 00
63 82 07 02 13 04 00 00 13 07 10 00 6F F0 5F F0
37 04 40 00 13 07 F0 0F 13 09 00 00 6F F0 5F EF
13 04 00 00 13 07 00 00 6F F0 9F EE 13 01 01 FE
23 28 21 01 13 59 75 01 23 2A 91 00 23 26 31 01
23 24 41 01 93 14 95 00 23 2E 11 00 23 2C 81 00
23 22 51 01 13 79 F9 0F 13 8A 05 00 93 D4 94 00
93 59 F5 01 63 06 09 08 93 07 F0 0F 63 02 F9 0A
93 94 34 00 B7 07 00 04 B3 E4 F4 00 13 09 19 F8
93 0A 00 00 13 55 7A 01 13 14 9A 00 13 75 F5 0F
13 54 94 00 13 5A FA 01 63 0C 05 08 93 07 F0 0F
63 08 F5 0A 13 14 34 00 B7 07 00 04 33 64 F4 00
13 05 15 F8 93 07 00 00 13 97 2A 00 33 67 F7 00
33 09 A9 00 13 07 F7 FF 93 06 E0 00 33 C8 49 01
93 08 19 00 63 EE E6 08 B7 16 40 00 13 17 27 00
93 86 46 84 33 07 D7 00 03 27 07 00 67 00 07 00
63 8A 04 02 13 85 04 00 EF 00 C0 33 93 07 B5 FF
13 09 A0 F8 B3 94 F4 00 33 09 A9 40 6F F0 5F F7
13 09 F0 0F 93 0A 20 00 E3 86 04 F6 93 0A 30 00
6F F0 5F F6 13 09 00 00 93 0A 10 00 6F F0 9F F5
63 0A 04 02 13 05 04 00 EF 00 C0 2F 93 07 B5 FF
33 14 F4 00 93 07 A0 F8 33 85 A7 40 6F F0 9F F6
13 05 F0 0F 93 07 20 00 E3 00 04 F6 93 07 30 00
6F F0 9F F5 13 05 00 00 93 07 10 00 6F F0 DF F4
37 0F 01 00 93 0E FF FF 93 DF 04 01 93 57 04 01
B3 F4 D4 01 33 74 D4 01 13 85 04 00 93 05 04 00
EF 00 C0 1C 13 03 05 00 93 85 07 00 13 85 04 00
EF 00 C0 1B 13 0E 05 00 93 05 04 00 13 85 0F 00
EF 00 C0 1A 13 07 05 00 93 85 07 00 13 85 0F 00
EF 00 C0 19 93 57 03 01 33 0E EE 00 B3 87 C7 01
63 F4 E7 00 33 05 E5 01 33 F7 D7 01 13 17 07 01
33 73 D3 01 33 07 67 00 13 14 67 00 33 34 80 00
93 D7 07 01 13 57 A7 01 33 67 E4 00 33 84 A7 00
13 14 64 00 33 64 E4 00 B7 07 00 08 B3 77 F4 00
63 8E 07 08 93 57 14 00 13 74 14 00 33 E4 87 00
13 87 F8 07 63 58 E0 08 93 77 74 00 63 8A 07 00
93 77 F4 00 93 06 40 00 63 84 D7 00 13 04 44 00
B7 07 00 08 B3 77 F4 00 63 8A 07 00 B7 07 00 F8
93 87 F7 FF 33 74 F4 00 13 87 08 08 93 07 E0 0F
13 54 34 00 63 DA E7 0A 13 04 00 00 13 07 F0 0F
6F 00 80 0A 13 88 09 00 13 84 04 00 93 87 0A 00
13 07 20 00 E3 82 E7 FE 13 07 30 00 63 80 E7 08
13 07 10 00 E3 96 E7 F8 13 04 00 00 13 07 00 00
6F 00 80 07 13 08 0A 00 6F F0 9F FD 93 08 09 00
6F F0 1F F7 93 07 10 00 B3 87 E7 40 13 07 B0 01
E3 4C F7 FC 93 88 E8 09 B3 57 F4 00 33 14 14 01
33 34 80 00 33 E4 87 00 93 77 74 00 63 8A 07 00
93 77 F4 00 13 07 40 00 63 84 E7 00 13 04 44 00
B7 07 00 04 B3 77 F4 00 13 54 34 00 E3 80 07 FA
13 04 00 00 13 07 10 00 6F 00 00 01 37 04 40 00
13 07 F0 0F 13 08 00 00 93 17 77 01 13 14 94 00
37 07 80 7F B3 F7 E7 00 13 54 94 00 33 E4 87 00
13 15 F8 01 83 20 C1 01 33 65 A4 00 03 24 81 01
83 24 41 01 03 29 01 01 83 29 C1 00 03 2A 81 00
83 2A 41 00 13 01 01 02 67 80 00 00 13 06 05 00
13 05 00 00 93 F6 15 00 63 84 06 00 33 05 C5 00
93 D5 15 00 13 16 16 00 E3 96 05 FE 67 80 00 00
63 40 05 06 63 C6 05 06 13 86 05 00 93 05 05 00
13 05 F0 FF 63 0C 06 02 93 06 10 00 63 7A B6 00
63 58 C0 00 13 16 16 00 93 96 16 00 E3 6A B6 FE
13 05 00 00 63 E6 C5 00 B3 85 C5 40 33 65 D5 00
93 D6 16 00 13 56 16 00 E3 96 06 FE 67 80 00 00
93 82 00 00 EF F0 5F FB 13 85 05 00 67 80 02 00
33 05 A0 40 63 48 B0 00 B3 05 B0 40 6F F0 DF F9
B3 05 B0 40 93 82 00 00 EF F0 1F F9 33 05 A0 40
67 80 02 00 93 82 00 00 63 CA 05 00 63 4C 05 00
EF F0 9F F7 13 85 05 00 67 80 02 00 B3 05 B0 40
E3 58 05 FE 33 05 A0 40 EF F0 1F F6 33 05 B0 40
67 80 02 00 B7 07 01 00 63 7A F5 02 93 07 F0 0F
B3 B7 A7 00 93 97 37 00 37 17 40 00 93 06 00 02
B3 86 F6 40 33 55 F5 00 93 07 07 88 33 85 A7 00
03 45 05 00 33 85 A6 40 67 80 00 00 37 07 00 01
93 07 00 01 E3 6A E5 FC 93 07 80 01 6F F0 DF FC
@00400800
00 00 C0 3F CD CC 0C 40 BC 08 00 00 48 09 00 00
C8 08 00 00 48 09 00 00 38 09 00 00 48 09 00 00
C8 08 00 00 BC 08 00 00 BC 08 00 00 38 09 00 00
C8 08 00 00 98 08 00 00 98 08 00 00 98 08 00 00
D0 08 00 00 A8 0B 00 00 A8 0B 00 00 CC 0B 00 00
A0 0B 00 00 A0 0B 00 00 34 0C 00 00 CC 0B 00 00
A0 0B 00 00 34 0C 00 00 A0 0B 00 00 CC 0B 00 00
9C 0B 00 00 9C 0B 00 00 9C 0B 00 00 34 0C 00 00
00 01 02 02 03 03 03 03 04 04 04 04 04 04 04 04
05 05 05 05 05 05 05 05 05 05 05 05 05 05 05 05
06 06 06 06 06 06 06 06 06 06 06 06 06 06 06 06
06 06 06 06 06 06 06 06 06 06 06 06 06 06 06 06
07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07
07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07
07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07
07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
