/*
 this module wrapps the UART IP 
 design and compacts the use of 
 uart via interface connections
 */

`timescale 1ns/1ns

module uart_wrapper
  #()
   (
    // slave wishbone interface
    // uart RX/TX signals
    );   
   
endmodule // uart_wrapper
