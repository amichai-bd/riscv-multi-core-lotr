//-----------------------------------------------------------------------------
// Title            : ring_controler 
// Project          : LOTR
//-----------------------------------------------------------------------------
// File             : ring_controler 
// Original Author  : Tzahi Peretz, Shimi Haleluya 
// Created          : 4/2021
//-----------------------------------------------------------------------------
// Description :
// The "ring_controler" implements :
// 
//------------------------------------------------------------------------------
// Modification history :
//
//
//------------------------------------------------------------------------------

module ring_controler 



endmodule
