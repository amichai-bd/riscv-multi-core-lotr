@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 00 0D 67 80 00 00
@0000001C
13 01 01 FE 23 2E 11 00 23 2C 81 00 23 2A 91 00
13 04 01 02 23 26 A4 FE 83 27 C4 FE 63 96 07 00
93 07 10 00 6F 00 40 04 03 27 C4 FE 93 07 10 00
63 16 F7 00 93 07 10 00 6F 00 00 03 83 27 C4 FE
93 87 F7 FF 13 85 07 00 EF F0 9F FB 93 04 05 00
83 27 C4 FE 93 87 E7 FF 13 85 07 00 EF F0 5F FA
93 07 05 00 B3 87 F4 00 13 85 07 00 83 20 C1 01
03 24 81 01 83 24 41 01 13 01 01 02 67 80 00 00
13 01 01 FE 23 2E 11 00 23 2C 81 00 13 04 01 02
13 05 60 00 EF F0 DF F6 93 07 05 00 23 26 F4 FE
B7 17 40 00 93 87 87 FF 03 27 C4 FE 23 A0 E7 00
93 07 00 00 13 85 07 00 83 20 C1 01 03 24 81 01
13 01 01 02 67 80 00 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 17 01 40 00 13 01 01 0E EF F0 5F F7
