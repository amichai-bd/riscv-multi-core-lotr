@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 50 68 73 00 10 00
@000000A8
13 01 01 FD 23 26 81 02 13 04 01 03 93 07 05 00
23 2C B4 FC 23 2A C4 FC A3 0F F4 FC 03 27 84 FD
93 07 07 00 93 97 27 00 B3 87 E7 00 93 97 67 00
23 26 F4 FE 83 27 44 FD 93 97 27 00 23 24 F4 FE
03 27 84 FE 83 27 C4 FE 33 07 F7 00 B7 07 40 03
B3 07 F7 00 23 22 F4 FE 03 27 84 FE 83 27 C4 FE
33 07 F7 00 B7 07 40 03 93 87 07 14 B3 07 F7 00
23 20 F4 FE 83 47 F4 FD 37 07 40 00 13 07 07 55
93 97 27 00 B3 07 F7 00 83 A7 07 00 13 87 07 00
83 27 44 FE 23 A0 E7 00 83 47 F4 FD 37 07 40 00
13 07 47 6D 93 97 27 00 B3 07 F7 00 83 A7 07 00
13 87 07 00 83 27 04 FE 23 A0 E7 00 13 00 00 00
03 24 C1 02 13 01 01 03 67 80 00 00 13 01 01 FD
23 26 11 02 23 24 81 02 13 04 01 03 23 2E A4 FC
23 26 04 FE 23 24 04 FE 23 22 04 FE B7 07 C0 00
93 87 07 22 83 A7 07 00 23 22 F4 FE B7 07 C0 00
93 87 47 23 83 A7 07 00 23 24 F4 FE 6F 00 80 0B
83 27 C4 FE 03 27 C4 FD B3 07 F7 00 03 C7 07 00
93 07 A0 00 63 1A F7 02 23 22 04 FE 83 27 84 FE
93 87 27 00 23 24 F4 FE 03 27 84 FE 93 07 80 07
63 14 F7 00 23 24 04 FE 83 27 C4 FE 93 87 17 00
23 26 F4 FE 6F 00 00 07 83 27 C4 FE 03 27 C4 FD
B3 07 F7 00 83 C7 07 00 03 27 84 FE 83 26 44 FE
13 86 06 00 93 05 07 00 13 85 07 00 EF F0 5F E8
83 27 44 FE 93 87 17 00 23 22 F4 FE 03 27 44 FE
93 07 00 05 63 12 F7 02 23 22 04 FE 83 27 84 FE
93 87 27 00 23 24 F4 FE 03 27 84 FE 93 07 80 07
63 14 F7 00 23 24 04 FE 83 27 C4 FE 93 87 17 00
23 26 F4 FE 83 27 C4 FE 03 27 C4 FD B3 07 F7 00
83 C7 07 00 E3 9E 07 F2 B7 07 C0 00 93 87 07 22
03 27 44 FE 23 A0 E7 00 B7 07 C0 00 93 87 47 23
03 27 84 FE 23 A0 E7 00 13 00 00 00 83 20 C1 02
03 24 81 02 13 01 01 03 67 80 00 00 13 01 01 FD
23 26 81 02 13 04 01 03 23 2E A4 FC 23 2C B4 FC
23 2A C4 FC 03 27 84 FD 93 07 07 00 93 97 27 00
B3 87 E7 00 93 97 67 00 23 26 F4 FE 83 27 44 FD
93 97 27 00 23 24 F4 FE 03 27 84 FE 83 27 C4 FE
33 07 F7 00 B7 07 40 03 B3 07 F7 00 23 22 F4 FE
03 27 84 FE 83 27 C4 FE 33 07 F7 00 B7 07 40 03
93 87 07 14 B3 07 F7 00 23 20 F4 FE B7 17 40 00
13 87 87 85 83 27 C4 FD 93 97 27 00 B3 07 F7 00
83 A7 07 00 13 87 07 00 83 27 44 FE 23 A0 E7 00
B7 17 40 00 13 87 07 87 83 27 C4 FD 93 97 27 00
B3 07 F7 00 83 A7 07 00 13 87 07 00 83 27 04 FE
23 A0 E7 00 13 00 00 00 03 24 C1 02 13 01 01 03
67 80 00 00 13 01 01 FE 23 2E 81 00 13 04 01 02
23 26 A4 FE 23 24 B4 FE B7 07 C0 00 93 87 07 22
03 27 84 FE 23 A0 E7 00 B7 07 C0 00 93 87 47 23
03 27 C4 FE 23 A0 E7 00 13 00 00 00 03 24 C1 01
13 01 01 02 67 80 00 00 13 01 01 FE 23 2E 81 00
13 04 01 02 23 26 04 FE B7 07 40 03 23 24 F4 FE
23 26 04 FE 6F 00 40 02 83 27 C4 FE 93 97 27 00
03 27 84 FE B3 07 F7 00 23 A0 07 00 83 27 C4 FE
93 87 17 00 23 26 F4 FE 03 27 C4 FE B7 27 00 00
93 87 F7 57 E3 DA E7 FC 13 00 00 00 13 00 00 00
03 24 C1 01 13 01 01 02 67 80 00 00 13 01 01 FC
23 2E 11 02 23 2C 81 02 13 04 01 04 23 26 A4 FC
23 26 04 FE 23 24 04 FE 83 27 C4 FC 63 D6 07 02
83 27 C4 FE 13 87 17 00 23 26 E4 FE 13 07 04 FF
B3 07 F7 00 13 07 D0 02 23 80 E7 FE 83 27 C4 FC
B3 07 F0 40 23 26 F4 FC 83 27 C4 FC 93 05 A0 00
13 85 07 00 EF 10 00 58 93 07 05 00 13 F7 F7 0F
83 27 C4 FE 93 86 17 00 23 26 D4 FE 13 07 07 03
13 77 F7 0F 93 06 04 FF B3 87 F6 00 23 80 E7 FE
83 27 C4 FC 93 05 A0 00 13 85 07 00 EF 10 40 4C
93 07 05 00 23 26 F4 FC 83 27 C4 FC E3 46 F0 FA
23 24 04 FE 6F 00 00 07 83 27 84 FE 13 07 04 FF
B3 07 F7 00 83 C7 07 FE A3 0F F4 FC 03 27 C4 FE
83 27 84 FE B3 07 F7 40 93 87 F7 FF 13 07 04 FF
B3 07 F7 00 03 C7 07 FE 83 27 84 FE 93 06 04 FF
B3 87 F6 00 23 80 E7 FE 03 27 C4 FE 83 27 84 FE
B3 07 F7 40 93 87 F7 FF 13 07 04 FF B3 07 F7 00
03 47 F4 FD 23 80 E7 FE 83 27 84 FE 93 87 17 00
23 24 F4 FE 83 27 C4 FE 13 D7 F7 01 B3 07 F7 00
93 D7 17 40 13 87 07 00 83 27 84 FE E3 CE E7 F6
B7 07 C0 00 93 87 47 23 83 A7 07 00 23 22 F4 FE
B7 07 C0 00 93 87 07 22 83 A7 07 00 23 20 F4 FE
23 24 04 FE 6F 00 80 06 83 27 84 FE 13 07 04 FF
B3 07 F7 00 83 C7 07 FE 03 26 04 FE 83 25 44 FE
13 85 07 00 EF F0 DF B0 83 27 04 FE 93 87 17 00
23 20 F4 FE 03 27 04 FE 93 07 00 05 63 1A F7 00
23 20 04 FE 83 27 44 FE 93 87 27 00 23 22 F4 FE
03 27 44 FE 93 07 70 07 63 D4 E7 00 23 22 04 FE
83 27 84 FE 93 87 17 00 23 24 F4 FE 03 27 84 FE
83 27 C4 FE E3 4A F7 F8 B7 07 C0 00 93 87 07 22
03 27 04 FE 23 A0 E7 00 B7 07 C0 00 93 87 47 23
03 27 44 FE 23 A0 E7 00 13 00 00 00 83 20 C1 03
03 24 81 03 13 01 01 04 67 80 00 00 13 01 01 FE
23 2E 81 00 13 04 01 02 23 26 04 FE 6F 00 00 01
83 27 C4 FE 93 87 17 00 23 26 F4 FE 03 27 C4 FE
B7 47 01 00 93 87 F7 87 E3 D4 E7 FE 13 00 00 00
13 00 00 00 03 24 C1 01 13 01 01 02 67 80 00 00
13 01 01 FD 23 26 81 02 13 04 01 03 23 2E A4 FC
23 2C B4 FC 23 2A C4 FC 23 28 D4 FC 83 27 84 FD
93 87 17 14 93 97 17 00 03 27 44 FD B3 07 F7 00
23 22 F4 FE 03 27 C4 FD 93 07 07 00 93 97 27 00
B3 87 E7 00 93 97 47 00 93 87 17 00 23 20 F4 FE
23 26 04 FE 6F 00 40 03 03 27 44 FE 83 27 C4 FE
33 07 F7 40 83 27 04 FD B3 07 F7 00 13 97 27 00
B7 07 40 03 B3 07 F7 00 23 A0 07 00 83 27 C4 FE
93 87 07 05 23 26 F4 FE 03 27 C4 FE 93 07 00 64
E3 D4 E7 FC 23 24 04 FE 6F 00 80 03 03 27 44 FE
83 27 84 FE 33 07 F7 40 83 27 04 FD B3 07 F7 00
13 97 27 00 B7 07 40 03 B3 07 F7 00 13 07 F0 FF
23 A0 E7 00 83 27 84 FE 93 87 07 05 23 24 F4 FE
03 27 84 FE 83 27 04 FE E3 42 F7 FC 13 00 00 00
13 00 00 00 03 24 C1 02 13 01 01 03 67 80 00 00
13 01 01 FD 23 26 81 02 13 04 01 03 23 2E A4 FC
23 2C B4 FC 83 27 C4 FD 83 A7 07 00 23 26 F4 FE
83 27 84 FD 03 A7 07 00 83 27 C4 FD 23 A0 E7 00
83 27 84 FD 03 27 C4 FE 23 A0 E7 00 13 00 00 00
03 24 C1 02 13 01 01 03 67 80 00 00 13 01 01 FD
23 26 11 02 23 24 81 02 13 04 01 03 23 2E A4 FC
23 2C B4 FC 23 2A C4 FC 23 28 D4 FC 23 26 04 FE
6F 00 C0 0F 23 24 04 FE 6F 00 00 0D 83 27 84 FE
93 97 27 00 03 27 C4 FD B3 07 F7 00 03 A7 07 00
83 27 84 FE 93 87 17 00 93 97 27 00 83 26 C4 FD
B3 87 F6 00 83 A7 07 00 63 DA E7 08 83 27 84 FE
93 97 27 00 03 27 C4 FD B3 06 F7 00 83 27 84 FE
93 87 17 00 93 97 27 00 03 27 C4 FD B3 07 F7 00
93 85 07 00 13 85 06 00 EF F0 9F F2 83 27 84 FE
93 97 27 00 03 27 C4 FD B3 07 F7 00 83 A7 07 00
83 26 04 FD 03 26 44 FD 83 25 84 FE 13 85 07 00
EF F0 1F E1 83 27 84 FE 93 87 17 00 93 97 27 00
03 27 C4 FD B3 07 F7 00 03 A7 07 00 83 27 84 FE
93 87 17 00 83 26 04 FD 03 26 44 FD 93 85 07 00
13 05 07 00 EF F0 DF DD EF F0 5F D9 83 27 84 FE
93 87 17 00 23 24 F4 FE 03 27 84 FD 83 27 C4 FE
B3 07 F7 40 93 87 F7 FF 03 27 84 FE E3 40 F7 F2
83 27 C4 FE 93 87 17 00 23 26 F4 FE 83 27 84 FD
93 87 F7 FF 03 27 C4 FE E3 4E F7 EE 13 00 00 00
13 00 00 00 83 20 C1 02 03 24 81 02 13 01 01 03
67 80 00 00 13 01 01 FD 23 26 11 02 23 24 81 02
13 04 01 03 23 2E A4 FC 23 2C B4 FC 23 2A C4 FC
23 28 D4 FC 93 07 10 00 23 26 F4 FE 6F 00 00 12
83 27 C4 FE 93 97 27 00 03 27 C4 FD B3 07 F7 00
83 A7 07 00 23 22 F4 FE 83 27 C4 FE 93 87 F7 FF
23 24 F4 FE 6F 00 40 07 83 27 84 FE 93 97 27 00
03 27 C4 FD 33 07 F7 00 83 27 84 FE 93 87 17 00
93 97 27 00 83 26 C4 FD B3 87 F6 00 03 27 07 00
23 A0 E7 00 83 27 84 FE 93 87 17 00 93 97 27 00
03 27 C4 FD B3 07 F7 00 03 A7 07 00 83 27 84 FE
93 87 17 00 83 26 04 FD 03 26 44 FD 93 85 07 00
13 05 07 00 EF F0 DF CC EF F0 5F C8 83 27 84 FE
93 87 F7 FF 23 24 F4 FE 83 27 84 FE 63 C0 07 02
83 27 84 FE 93 97 27 00 03 27 C4 FD B3 07 F7 00
83 A7 07 00 03 27 44 FE E3 48 F7 F6 83 27 84 FE
93 87 17 00 93 97 27 00 03 27 C4 FD B3 07 F7 00
03 27 44 FE 23 A0 E7 00 83 27 84 FE 93 87 17 00
93 97 27 00 03 27 C4 FD B3 07 F7 00 03 A7 07 00
83 27 84 FE 93 87 17 00 83 26 04 FD 03 26 44 FD
93 85 07 00 13 05 07 00 EF F0 9F C4 EF F0 1F C0
83 27 C4 FE 93 87 17 00 23 26 F4 FE 03 27 C4 FE
83 27 84 FD E3 4E F7 EC 13 00 00 00 13 00 00 00
83 20 C1 02 03 24 81 02 13 01 01 03 67 80 00 00
13 01 01 FF 23 26 11 00 23 24 81 00 13 04 01 01
93 05 10 00 13 05 10 00 EF F0 DF 90 B7 07 40 00
13 85 07 00 EF F0 8F EF 93 05 10 00 13 05 A0 00
EF F0 5F 8F B7 07 40 00 13 85 C7 01 EF F0 0F EE
93 05 40 01 13 05 40 01 EF F0 DF 8D B7 07 40 00
13 85 C7 03 EF F0 8F EC 93 05 40 01 13 05 80 02
EF F0 5F 8C B7 07 40 00 13 85 C7 05 EF F0 0F EB
93 05 40 01 13 05 20 03 EF F0 DF 8A B7 07 40 00
13 85 87 07 EF F0 8F E9 93 05 40 01 13 05 C0 03
EF F0 5F 89 B7 07 40 00 13 85 87 08 EF F0 0F E8
93 05 40 01 13 05 60 04 EF F0 DF 87 B7 07 40 00
13 85 07 0A EF F0 8F E6 13 00 00 00 83 20 C1 00
03 24 81 00 13 01 01 01 67 80 00 00 13 01 01 FD
23 26 11 02 23 24 81 02 13 04 01 03 93 07 10 00
23 26 F4 FE 93 07 F0 3F 23 24 F4 FE 23 22 04 FE
93 07 10 00 23 20 F4 FE 93 07 00 20 23 2E F4 FC
93 05 A0 00 13 05 40 01 EF F0 DF 81 B7 07 40 00
13 85 47 0B EF F0 8F E0 93 05 F0 00 13 05 E0 01
EF F0 5F 80 B7 07 40 00 13 85 07 0D EF F0 0F DF
93 05 40 01 13 05 80 02 EF F0 CF FE B7 07 40 00
13 85 47 10 EF F0 8F DD 93 05 40 01 13 05 D0 02
EF F0 4F FD B7 07 40 00 13 85 C7 11 EF F0 0F DC
93 05 40 01 13 05 20 03 EF F0 CF FB B7 07 40 00
13 85 47 13 EF F0 8F DA 93 05 40 01 13 05 70 03
EF F0 4F FA B7 07 40 00 13 85 07 15 EF F0 0F D9
B7 27 C0 03 93 87 47 02 83 A7 07 00 63 9C 07 04
93 07 10 00 23 26 F4 FE 93 07 F0 3F 23 24 F4 FE
93 07 10 00 23 20 F4 FE 93 07 00 20 23 2E F4 FC
EF F0 DF A0 B7 27 C0 03 93 87 87 01 03 27 44 FE
23 A0 E7 00 03 27 44 FE 93 07 F0 3F 63 16 F7 00
23 22 04 FE 6F F0 DF FA 93 07 F0 3F 23 22 F4 FE
6F F0 1F FA B7 27 C0 03 93 87 47 02 03 A7 07 00
93 07 10 00 63 1C F7 04 93 07 F0 3F 23 24 F4 FE
23 22 04 FE 93 07 10 00 23 20 F4 FE 93 07 00 20
23 2E F4 FC EF F0 9F 9A B7 27 C0 03 93 87 87 01
03 27 C4 FE 23 A0 E7 00 83 27 C4 FE 93 87 17 00
23 26 F4 FE 03 27 C4 FE 93 07 F0 3F E3 12 F7 F4
93 07 10 00 23 26 F4 FE 6F F0 9F F3 B7 27 C0 03
93 87 47 02 03 A7 07 00 93 07 20 00 63 1C F7 04
93 07 10 00 23 26 F4 FE 93 07 F0 3F 23 24 F4 FE
23 22 04 FE 93 07 00 20 23 2E F4 FC EF F0 1F 94
B7 27 C0 03 93 87 87 01 03 27 04 FE 23 A0 E7 00
83 27 04 FE 93 97 17 00 23 20 F4 FE 03 27 04 FE
93 07 00 20 E3 DE E7 EC 93 07 10 00 23 20 F4 FE
6F F0 1F ED B7 27 C0 03 93 87 47 02 03 A7 07 00
93 07 30 00 E3 1E F7 EA 93 07 10 00 23 26 F4 FE
23 22 04 FE 93 07 10 00 23 20 F4 FE 93 07 00 20
23 2E F4 FC EF F0 9F 8D B7 27 C0 03 93 87 87 01
03 27 84 FE 23 A0 E7 00 83 27 84 FE 93 87 F7 FF
23 24 F4 FE 83 27 84 FE E3 9C 07 E6 93 07 F0 3F
23 24 F4 FE 6F F0 DF E6 13 01 01 FF 23 26 11 00
23 24 81 00 13 04 01 01 93 05 10 00 13 05 10 00
EF F0 4F DE B7 07 40 00 13 85 07 17 EF F0 0F BD
93 05 10 00 13 05 50 00 EF F0 CF DC B7 07 40 00
13 85 07 18 EF F0 8F BB 93 05 40 01 13 05 A0 00
EF F0 4F DB B7 07 40 00 13 85 87 18 EF F0 0F BA
93 05 40 01 13 05 40 01 EF F0 CF D9 B7 07 40 00
13 85 07 1A EF F0 8F B8 93 05 40 01 13 05 90 01
EF F0 4F D8 B7 07 40 00 13 85 47 1B EF F0 0F B7
93 05 40 01 13 05 E0 01 EF F0 CF D6 B7 07 40 00
13 85 47 1D EF F0 8F B5 93 05 40 01 13 05 30 02
EF F0 4F D5 B7 07 40 00 13 85 C7 1E EF F0 0F B4
93 05 40 01 13 05 80 02 EF F0 CF D3 B7 07 40 00
13 85 C7 21 EF F0 8F B2 93 05 40 01 13 05 D0 02
EF F0 4F D2 B7 07 40 00 13 85 47 24 EF F0 0F B1
93 05 40 01 13 05 20 03 EF F0 CF D0 B7 07 40 00
13 85 07 26 EF F0 8F AF 93 05 90 01 13 05 70 03
EF F0 4F CF B7 07 40 00 13 85 87 27 EF F0 0F AE
93 05 90 01 13 05 C0 03 EF F0 CF CD B7 07 40 00
13 85 C7 28 EF F0 8F AC 93 05 40 01 13 05 10 04
EF F0 4F CC B7 07 40 00 13 85 07 2A EF F0 0F AB
93 05 90 01 13 05 60 04 EF F0 CF CA B7 07 40 00
13 85 C7 2A EF F0 8F A9 93 05 90 01 13 05 B0 04
EF F0 4F C9 B7 07 40 00 13 85 87 2B EF F0 0F A8
93 05 90 01 13 05 00 05 EF F0 CF C7 B7 07 40 00
13 85 87 2C EF F0 8F A6 13 00 00 00 83 20 C1 00
03 24 81 00 13 01 01 01 67 80 00 00 13 01 01 F7
23 26 11 08 23 24 81 08 13 04 01 09 EF F0 CF C8
B7 07 C0 00 83 A7 07 00 23 24 F4 FC 93 07 20 01
23 22 F4 FC 83 27 84 FC 93 87 C7 FF 13 07 70 00
E3 60 F7 20 13 97 27 00 B7 07 40 00 93 87 07 53
B3 07 F7 00 83 A7 07 00 67 80 07 00 B7 07 C0 01
93 87 07 15 23 A0 07 00 EF F0 4F EA 93 05 10 00
13 05 E0 01 EF F0 0F BF B7 07 40 00 13 85 C7 2D
EF F0 CF 9D B7 07 40 00 13 87 07 41 93 07 84 F7
93 06 07 00 13 07 80 04 13 06 07 00 93 85 06 00
13 85 07 00 EF 00 10 27 23 24 04 FE 6F 00 C0 03
83 27 84 FE 93 97 27 00 13 07 04 FF B3 07 F7 00
03 A7 87 F8 B7 17 00 00 93 86 07 E1 13 06 00 00
83 25 84 FE 13 05 07 00 EF F0 8F E7 83 27 84 FE
93 87 17 00 23 24 F4 FE 03 27 84 FE 83 27 44 FC
E3 40 F7 FC EF F0 8F E1 13 07 84 F7 B7 17 00 00
93 86 07 E1 13 06 00 00 83 25 44 FC 13 05 07 00
EF F0 CF F7 EF F0 8F DF 6F 00 00 00 EF F0 5F A2
23 20 04 FC B7 27 C0 03 93 87 47 02 83 A7 07 00
23 20 F4 FC 03 27 04 FC 93 07 10 00 63 14 F7 04
13 06 20 01 93 05 80 02 13 05 10 00 EF F0 0F A5
13 06 20 01 93 05 20 03 13 05 50 00 EF F0 0F A4
13 06 20 01 93 05 C0 03 13 05 50 00 EF F0 0F A3
13 06 20 01 93 05 60 04 13 05 50 00 EF F0 0F A2
6F F0 5F FA 03 27 04 FC 93 07 20 00 63 14 F7 04
13 06 20 01 93 05 20 03 13 05 10 00 EF F0 0F A0
13 06 20 01 93 05 80 02 13 05 50 00 EF F0 0F 9F
13 06 20 01 93 05 C0 03 13 05 50 00 EF F0 0F 9E
13 06 20 01 93 05 60 04 13 05 50 00 EF F0 0F 9D
6F F0 5F F5 03 27 04 FC 93 07 40 00 63 14 F7 04
13 06 20 01 93 05 C0 03 13 05 10 00 EF F0 0F 9B
13 06 20 01 93 05 80 02 13 05 50 00 EF F0 0F 9A
13 06 20 01 93 05 20 03 13 05 50 00 EF F0 0F 99
13 06 20 01 93 05 60 04 13 05 50 00 EF F0 0F 98
6F F0 5F F0 03 27 04 FC 93 07 50 00 63 14 F7 04
13 06 20 01 93 05 60 04 13 05 10 00 EF F0 0F 96
13 06 20 01 93 05 80 02 13 05 50 00 EF F0 0F 95
13 06 20 01 93 05 20 03 13 05 50 00 EF F0 0F 94
13 06 20 01 93 05 C0 03 13 05 50 00 EF F0 0F 93
6F F0 5F EB 03 27 04 FC 93 07 10 08 63 06 F7 06
03 27 04 FC 93 07 20 08 63 00 F7 06 03 27 04 FC
93 07 40 08 63 0A F7 04 03 27 04 FC 93 07 50 08
63 04 F7 04 13 06 20 01 93 05 80 02 13 05 50 00
EF F0 CF 8E 13 06 20 01 93 05 20 03 13 05 50 00
EF F0 CF 8D 13 06 20 01 93 05 C0 03 13 05 50 00
EF F0 CF 8C 13 06 20 01 93 05 60 04 13 05 50 00
EF F0 CF 8B 6F F0 1F E4 03 27 04 FC 93 07 10 08
63 18 F7 00 EF F0 4F 9B EF F0 1F B7 6F 00 00 00
03 27 04 FC 93 07 20 08 63 18 F7 00 EF F0 CF 99
EF F0 DF 8F 6F 00 00 00 03 27 04 FC 93 07 50 08
63 1C F7 00 EF F0 4F 98 B7 07 40 00 13 85 87 2F
EF E0 DF F2 6F 00 00 00 03 27 04 FC 93 07 40 08
63 12 F7 70 EF F0 4F 96 B7 07 C0 02 13 87 C7 15
93 07 10 00 23 20 F7 00 37 07 C0 02 13 07 87 15
23 20 F7 00 37 07 C0 02 13 07 47 15 23 20 F7 00
37 07 C0 02 13 07 07 15 23 20 F7 00 37 07 C0 01
13 07 C7 15 23 20 F7 00 37 07 C0 01 13 07 87 15
23 20 F7 00 37 07 C0 01 13 07 07 15 23 20 F7 00
EF F0 CF B6 93 05 80 02 13 05 A0 05 EF F0 8F 8B
B7 07 40 00 13 85 87 32 EF E0 5F EA B7 07 40 00
13 87 87 45 93 07 84 F7 93 06 07 00 13 07 80 04
13 06 07 00 93 85 06 00 13 85 07 00 EF 00 80 73
23 22 04 FE 6F 00 00 04 83 27 44 FE 93 97 27 00
13 07 04 FF B3 07 F7 00 03 A7 87 F8 B7 17 00 00
93 86 07 E1 B7 17 00 00 13 86 87 2E 83 25 44 FE
13 05 07 00 EF F0 CF B3 83 27 44 FE 93 87 17 00
23 22 F4 FE 03 27 44 FE 83 27 44 FC E3 4E F7 FA
EF F0 CF AD 13 07 84 F7 B7 17 00 00 93 86 07 E1
B7 17 00 00 13 86 87 2E 83 25 44 FC 13 05 07 00
EF F0 CF C3 EF F0 8F AB 6F 00 00 00 B7 07 C0 01
93 87 87 15 23 A0 07 00 23 26 04 FE 6F 00 C0 0B
83 27 C4 FE 13 97 27 00 B7 07 40 03 B3 07 F7 00
13 07 F0 FF 23 A0 E7 00 03 27 C4 FE B7 17 00 00
93 87 07 96 B3 07 F7 00 13 97 27 00 B7 07 40 03
93 87 07 EC B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
03 27 C4 FE B7 17 00 00 93 87 07 2C B3 07 F7 00
13 97 27 00 B7 07 40 03 93 87 07 EC B3 07 F7 00
13 07 F0 FF 23 A0 E7 00 03 27 C4 FE B7 27 00 00
93 87 07 C2 B3 07 F7 00 13 97 27 00 B7 07 40 03
93 87 07 EC B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
83 27 C4 FE 13 97 27 00 B7 97 40 03 93 87 07 4C
B3 07 F7 00 13 07 F0 FF 23 A0 E7 00 83 27 C4 FE
93 87 17 00 23 26 F4 FE 03 27 C4 FE 93 07 F0 04
E3 D0 E7 F4 23 26 04 FE 6F 00 00 09 03 27 C4 FE
93 07 07 00 93 97 27 00 B3 87 E7 00 93 97 67 00
13 87 07 00 B7 07 40 03 B3 07 F7 00 13 07 F0 FF
23 A0 E7 00 03 27 C4 FE 93 07 07 00 93 97 27 00
B3 87 E7 00 93 97 67 00 13 87 07 00 B7 07 40 03
93 87 C7 09 B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
03 27 C4 FE 93 07 07 00 93 97 27 00 B3 87 E7 00
93 97 67 00 13 87 07 00 B7 07 40 03 93 87 C7 13
B3 07 F7 00 13 07 F0 FF 23 A0 E7 00 83 27 C4 FE
93 87 17 00 23 26 F4 FE 03 27 C4 FE 93 07 70 07
E3 D6 E7 F6 EF F0 8F 93 93 05 80 02 13 05 E0 01
EF E0 5F E8 B7 07 40 00 13 85 87 34 EF E0 1F C7
B7 07 40 00 13 87 07 4A 93 07 84 F7 93 06 07 00
13 07 80 04 13 06 07 00 93 85 06 00 13 85 07 00
EF 00 40 50 23 20 04 FE 6F 00 C0 03 83 27 04 FE
93 97 27 00 13 07 04 FF B3 07 F7 00 03 A7 87 F8
B7 17 00 00 93 86 07 E1 13 06 80 02 83 25 04 FE
13 05 07 00 EF F0 CF 90 83 27 04 FE 93 87 17 00
23 20 F4 FE 03 27 04 FE 83 27 44 FC E3 40 F7 FC
EF F0 CF 8A 13 07 84 F7 B7 17 00 00 93 86 07 E1
13 06 80 02 83 25 44 FC 13 05 07 00 EF F0 0F A1
EF F0 CF 88 6F 00 00 00 B7 07 C0 01 93 87 C7 15
23 A0 07 00 EF F0 8F 87 93 05 10 00 13 05 A0 05
EF E0 5F DC B7 07 40 00 13 85 47 36 EF E0 1F BB
B7 07 40 00 13 87 87 4E 93 07 84 F7 93 06 07 00
13 07 80 04 13 06 07 00 93 85 06 00 13 85 07 00
EF 00 40 44 23 2E 04 FC 6F 00 00 04 83 27 C4 FD
93 97 27 00 13 07 04 FF B3 07 F7 00 03 A7 87 F8
B7 17 00 00 93 86 07 E1 B7 17 00 00 13 86 07 2C
83 25 C4 FD 13 05 07 00 EF F0 8F 84 83 27 C4 FD
93 87 17 00 23 2E F4 FC 03 27 C4 FD 83 27 44 FC
E3 4E F7 FA EF E0 9F FE 13 07 84 F7 B7 17 00 00
93 86 07 E1 B7 17 00 00 13 86 07 2C 83 25 44 FC
13 05 07 00 EF F0 8F 94 EF E0 5F FC 6F 00 00 00
B7 07 C0 02 93 87 07 15 23 A0 07 00 EF E0 1F FB
93 05 10 00 13 05 10 00 EF E0 DF CF B7 07 40 00
13 85 87 38 EF E0 9F AE B7 07 40 00 13 87 07 41
93 07 84 F7 93 06 07 00 13 07 80 04 13 06 07 00
93 85 06 00 13 85 07 00 EF 00 C0 37 23 2C 04 FC
6F 00 80 03 83 27 84 FD 93 97 27 00 13 07 04 FF
B3 07 F7 00 83 A7 87 F8 93 06 00 4B 13 06 00 00
83 25 84 FD 13 85 07 00 EF E0 9F F8 83 27 84 FD
93 87 17 00 23 2C F4 FC 03 27 84 FD 83 27 44 FC
E3 42 F7 FC EF E0 9F F2 93 07 84 F7 93 06 00 4B
13 06 00 00 83 25 44 FC 13 85 07 00 EF F0 8F 9D
EF E0 DF F0 6F 00 00 00 B7 07 C0 02 93 87 47 15
23 A0 07 00 EF E0 9F EF 93 05 80 02 13 05 C0 03
EF E0 5F C4 B7 07 40 00 13 85 87 3A EF E0 1F A3
B7 07 40 00 13 87 87 45 93 07 84 F7 93 06 07 00
13 07 80 04 13 06 07 00 93 85 06 00 13 85 07 00
EF 00 40 2C 23 2A 04 FC 6F 00 C0 03 83 27 44 FD
93 97 27 00 13 07 04 FF B3 07 F7 00 03 A7 87 F8
93 06 00 4B B7 17 00 00 13 86 87 2E 83 25 44 FD
13 05 07 00 EF E0 DF EC 83 27 44 FD 93 87 17 00
23 2A F4 FC 03 27 44 FD 83 27 44 FC E3 40 F7 FC
EF E0 DF E6 13 07 84 F7 93 06 00 4B B7 17 00 00
13 86 87 2E 83 25 44 FC 13 05 07 00 EF F0 8F 91
EF E0 DF E4 6F 00 00 00 B7 07 C0 02 93 87 87 15
23 A0 07 00 EF E0 9F E3 93 05 80 02 13 05 10 00
EF E0 5F B8 B7 07 40 00 13 85 87 3C EF E0 1F 97
B7 07 40 00 13 87 07 4A 93 07 84 F7 93 06 07 00
13 07 80 04 13 06 07 00 93 85 06 00 13 85 07 00
EF 00 40 20 23 28 04 FC 6F 00 80 03 83 27 04 FD
93 97 27 00 13 07 04 FF B3 07 F7 00 83 A7 87 F8
93 06 00 4B 13 06 80 02 83 25 04 FD 13 85 07 00
EF E0 1F E1 83 27 04 FD 93 87 17 00 23 28 F4 FC
03 27 04 FD 83 27 44 FC E3 42 F7 FC EF E0 1F DB
93 07 84 F7 93 06 00 4B 13 06 80 02 83 25 44 FC
13 85 07 00 EF F0 0F 86 EF E0 5F D9 6F 00 00 00
B7 07 C0 02 93 87 C7 15 23 A0 07 00 EF E0 1F D8
93 05 10 00 13 05 C0 03 EF E0 DF AC B7 07 40 00
13 85 87 3E EF E0 9F 8B B7 07 40 00 13 87 87 4E
93 07 84 F7 93 06 07 00 13 07 80 04 13 06 07 00
93 85 06 00 13 85 07 00 EF 00 C0 14 23 26 04 FC
6F 00 C0 03 83 27 C4 FC 93 97 27 00 13 07 04 FF
B3 07 F7 00 03 A7 87 F8 93 06 00 4B B7 17 00 00
13 86 07 2C 83 25 C4 FC 13 05 07 00 EF E0 5F D5
83 27 C4 FC 93 87 17 00 23 26 F4 FC 03 27 C4 FC
83 27 44 FC E3 40 F7 FC EF E0 5F CF 13 07 84 F7
93 06 00 4B B7 17 00 00 13 86 07 2C 83 25 44 FC
13 05 07 00 EF E0 1F FA EF E0 5F CD 6F 00 00 00
6F 00 00 00 13 00 00 00 93 07 00 00 13 85 07 00
83 20 C1 08 03 24 81 08 13 01 01 09 67 80 00 00
63 40 05 06 63 C6 05 06 13 86 05 00 93 05 05 00
13 05 F0 FF 63 0C 06 02 93 06 10 00 63 7A B6 00
63 58 C0 00 13 16 16 00 93 96 16 00 E3 6A B6 FE
13 05 00 00 63 E6 C5 00 B3 85 C5 40 33 65 D5 00
93 D6 16 00 13 56 16 00 E3 96 06 FE 67 80 00 00
93 82 00 00 EF F0 5F FB 13 85 05 00 67 80 02 00
33 05 A0 40 63 48 B0 00 B3 05 B0 40 6F F0 DF F9
B3 05 B0 40 93 82 00 00 EF F0 1F F9 33 05 A0 40
67 80 02 00 93 82 00 00 63 CA 05 00 63 4C 05 00
EF F0 9F F7 13 85 05 00 67 80 02 00 B3 05 B0 40
E3 58 05 FE 33 05 A0 40 EF F0 1F F6 33 05 B0 40
67 80 02 00
@00001A2C
B3 C7 A5 00 93 F7 37 00 B3 08 C5 00 63 96 07 06
93 07 30 00 63 F2 C7 06 93 77 35 00 13 07 05 00
63 9A 07 0C 13 F6 C8 FF B3 06 E6 40 93 07 00 02
93 02 00 02 63 C2 D7 06 93 86 05 00 93 07 07 00
63 78 C7 02 03 A8 06 00 93 87 47 00 93 86 46 00
23 AE 07 FF E3 E8 C7 FE 93 07 F6 FF B3 87 E7 40
93 F7 C7 FF 93 87 47 00 33 07 F7 00 B3 85 F5 00
63 68 17 01 67 80 00 00 13 07 05 00 E3 7C 15 FF
83 C7 05 00 13 07 17 00 93 85 15 00 A3 0F F7 FE
E3 68 17 FF 67 80 00 00 83 A6 45 00 83 A7 C5 01
83 AF 05 00 03 AF 85 00 83 AE C5 00 03 AE 05 01
03 A3 45 01 03 A8 85 01 23 22 D7 00 83 A6 05 02
23 20 F7 01 23 24 E7 01 23 26 D7 01 23 28 C7 01
23 2A 67 00 23 2C 07 01 23 2E F7 00 13 07 47 02
B3 07 E6 40 23 2E D7 FE 93 85 45 02 E3 C6 F2 FA
6F F0 9F F4 83 C6 05 00 13 07 17 00 93 77 37 00
A3 0F D7 FE 93 85 15 00 E3 8E 07 F0 83 C6 05 00
13 07 17 00 93 77 37 00 A3 0F D7 FE 93 85 15 00
E3 9A 07 FC 6F F0 1F F0
