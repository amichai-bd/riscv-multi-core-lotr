@00000000
B7 07 00 00 93 87 07 00 63 8A 07 00 37 05 00 00
13 05 05 4A 17 03 00 00 67 00 43 47 67 80 00 00
97 21 00 00 93 81 81 DC 17 25 00 00 13 05 45 9F
17 26 00 00 13 06 86 A0 33 06 A6 40 93 05 00 00
97 00 00 00 E7 80 80 24 17 05 00 00 13 05 05 44
63 0A 05 00 17 05 00 00 13 05 C5 44 97 00 00 00
E7 80 C0 42 97 00 00 00 E7 80 80 18 03 25 01 00
93 05 41 00 13 06 00 00 97 00 00 00 E7 80 C0 08
17 03 00 00 67 00 03 13 B7 27 00 00 03 C7 C7 A1
63 14 07 04 13 01 01 FF 23 24 81 00 13 84 07 00
B7 07 00 00 23 26 11 00 93 87 07 00 63 8A 07 00
37 15 00 00 13 05 85 5D 97 00 00 00 E7 00 00 00
93 07 10 00 83 20 C1 00 23 0E F4 A0 03 24 81 00
13 01 01 01 67 80 00 00 67 80 00 00 B7 07 00 00
93 87 07 00 63 8E 07 00 B7 25 00 00 37 15 00 00
93 85 05 A2 13 05 85 5D 17 03 00 00 67 00 00 00
67 80 00 00 13 01 01 FE 23 2E 11 00 23 2C 81 00
13 04 01 02 93 07 50 00 23 26 F4 FE 93 07 30 00
23 24 F4 FE 83 25 84 FE 03 25 C4 FE 97 00 00 00
E7 80 00 06 93 07 05 00 23 22 F4 FE 93 07 50 00
23 26 F4 FE 93 07 30 00 23 24 F4 FE 83 25 84 FE
03 25 C4 FE 97 00 00 00 E7 80 80 03 93 07 05 00
23 22 F4 FE B7 17 00 00 93 87 07 F0 03 27 44 FE
23 A0 E7 00 93 07 00 00 13 85 07 00 83 20 C1 01
03 24 81 01 13 01 01 02 67 80 00 00 13 06 05 00
13 05 00 00 93 F6 15 00 63 84 06 00 33 05 C5 00
93 D5 15 00 13 16 16 00 E3 96 05 FE 67 80 00 00
13 01 01 FF 93 05 00 00 23 24 81 00 23 26 11 00
13 04 05 00 97 00 00 00 E7 80 00 1A B7 27 00 00
03 A5 07 A1 83 27 C5 03 63 84 07 00 E7 80 07 00
13 05 04 00 97 00 00 00 E7 80 40 3B 13 01 01 FF
23 24 81 00 23 20 21 01 37 14 00 00 37 19 00 00
93 07 C4 5D 13 09 C9 5D 33 09 F9 40 23 26 11 00
23 22 91 00 13 59 29 40 63 00 09 02 13 04 C4 5D
93 04 00 00 83 27 04 00 93 84 14 00 13 04 44 00
E7 80 07 00 E3 18 99 FE 37 14 00 00 37 19 00 00
93 07 C4 5D 13 09 49 5E 33 09 F9 40 13 59 29 40
63 00 09 02 13 04 C4 5D 93 04 00 00 83 27 04 00
93 84 14 00 13 04 44 00 E7 80 07 00 E3 18 99 FE
83 20 C1 00 03 24 81 00 83 24 41 00 03 29 01 00
13 01 01 01 67 80 00 00 13 03 F0 00 13 07 05 00
63 7E C3 02 93 77 F7 00 63 90 07 0A 63 92 05 08
93 76 06 FF 13 76 F6 00 B3 86 E6 00 23 20 B7 00
23 22 B7 00 23 24 B7 00 23 26 B7 00 13 07 07 01
E3 66 D7 FE 63 14 06 00 67 80 00 00 B3 06 C3 40
93 96 26 00 97 02 00 00 B3 86 56 00 67 80 C6 00
23 07 B7 00 A3 06 B7 00 23 06 B7 00 A3 05 B7 00
23 05 B7 00 A3 04 B7 00 23 04 B7 00 A3 03 B7 00
23 03 B7 00 A3 02 B7 00 23 02 B7 00 A3 01 B7 00
23 01 B7 00 A3 00 B7 00 23 00 B7 00 67 80 00 00
93 F5 F5 0F 93 96 85 00 B3 E5 D5 00 93 96 05 01
B3 E5 D5 00 6F F0 DF F6 93 96 27 00 97 02 00 00
B3 86 56 00 93 82 00 00 E7 80 06 FA 93 80 02 00
93 87 07 FF 33 07 F7 40 33 06 F6 00 E3 78 C3 F6
6F F0 DF F3 13 01 01 FD B7 27 00 00 23 2C 41 01
03 AA 07 A1 23 20 21 03 23 26 11 02 03 29 8A 14
23 24 81 02 23 22 91 02 23 2E 31 01 23 2A 51 01
23 28 61 01 23 26 71 01 23 24 81 01 63 00 09 04
13 0B 05 00 93 8B 05 00 93 0A 10 00 93 09 F0 FF
83 24 49 00 13 84 F4 FF 63 42 04 02 93 94 24 00
B3 04 99 00 63 84 0B 04 83 A7 44 10 63 80 77 05
13 04 F4 FF 93 84 C4 FF E3 16 34 FF 83 20 C1 02
03 24 81 02 83 24 41 02 03 29 01 02 83 29 C1 01
03 2A 81 01 83 2A 41 01 03 2B 01 01 83 2B C1 00
03 2C 81 00 13 01 01 03 67 80 00 00 83 27 49 00
83 A6 44 00 93 87 F7 FF 63 8E 87 04 23 A2 04 00
E3 88 06 FA 83 27 89 18 33 97 8A 00 03 2C 49 00
B3 77 F7 00 63 92 07 02 E7 80 06 00 03 27 49 00
83 27 8A 14 63 14 87 01 E3 84 27 F9 E3 88 07 F8
13 89 07 00 6F F0 DF F5 83 27 C9 18 83 A5 44 08
33 77 F7 00 63 1C 07 00 13 05 0B 00 E7 80 06 00
6F F0 DF FC 23 22 89 00 6F F0 9F FA 13 85 05 00
E7 80 06 00 6F F0 9F FB 93 05 05 00 93 06 00 00
13 06 00 00 13 05 00 00 17 03 00 00 67 00 43 06
13 01 01 FF 23 24 81 00 B7 17 00 00 37 14 00 00
13 04 44 5E 93 87 87 5E B3 87 87 40 23 22 91 00
23 26 11 00 93 D4 27 40 63 80 04 02 93 87 C7 FF
33 84 87 00 83 27 04 00 93 84 F4 FF 13 04 C4 FF
E7 80 07 00 E3 98 04 FE 83 20 C1 00 03 24 81 00
83 24 41 00 13 01 01 01 67 80 00 00 B7 27 00 00
03 A7 07 A1 83 27 87 14 63 8C 07 04 03 A7 47 00
13 08 F0 01 63 4E E8 06 13 18 27 00 63 06 05 02
33 83 07 01 23 24 C3 08 83 A8 87 18 13 06 10 00
33 16 E6 00 B3 E8 C8 00 23 A4 17 19 23 24 D3 10
93 06 20 00 63 04 D5 02 13 07 17 00 23 A2 E7 00
B3 87 07 01 23 A4 B7 00 13 05 00 00 67 80 00 00
93 07 C7 14 23 24 F7 14 6F F0 5F FA 83 A6 C7 18
13 07 17 00 23 A2 E7 00 33 E6 C6 00 23 A6 C7 18
B3 87 07 01 23 A4 B7 00 13 05 00 00 67 80 00 00
13 05 F0 FF 67 80 00 00 93 08 D0 05 73 00 00 00
63 44 05 00 6F 00 00 00 13 01 01 FF 23 24 81 00
13 04 05 00 23 26 11 00 33 04 80 40 97 00 00 00
E7 80 00 01 23 20 85 00 6F 00 00 00 B7 27 00 00
03 A5 87 A1 67 80 00 00
@000015D8
00 00 00 00
@000015DC
00 00 00 00 DC 00 00 00
@000015E4
88 00 00 00
@000015E8
00 00 00 00 D4 18 00 00 3C 19 00 00 A4 19 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 01 00 00 00 00 00 00 00
0E 33 CD AB 34 12 6D E6 EC DE 05 00 0B 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00
@00001A10
E8 15 00 00 00 00 00 00 E8 15 00 00
