@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 80 13 73 00 10 00
@000000A8
13 01 01 FE 23 2E 11 00 23 2C 81 00 13 04 01 02
93 07 40 01 23 26 F4 FE 93 07 50 00 23 24 F4 FE
83 25 84 FE 03 25 C4 FE EF 00 40 26 93 07 05 00
23 22 F4 FE 83 27 44 FE 13 85 07 00 83 20 C1 01
03 24 81 01 13 01 01 02 67 80 00 00 13 01 01 FE
23 2E 11 00 23 2C 81 00 13 04 01 02 93 07 80 00
23 26 F4 FE 93 07 90 01 23 24 F4 FE 83 25 84 FE
03 25 C4 FE EF 00 80 21 93 07 05 00 23 22 F4 FE
83 27 44 FE 13 85 07 00 83 20 C1 01 03 24 81 01
13 01 01 02 67 80 00 00 13 01 01 FE 23 2E 11 00
23 2C 81 00 13 04 01 02 93 07 A0 00 23 26 F4 FE
93 07 E0 01 23 24 F4 FE 83 25 84 FE 03 25 C4 FE
EF 00 C0 1C 93 07 05 00 23 22 F4 FE 83 27 44 FE
13 85 07 00 83 20 C1 01 03 24 81 01 13 01 01 02
67 80 00 00 13 01 01 FE 23 2E 11 00 23 2C 81 00
13 04 01 02 93 07 40 06 23 26 F4 FE 93 07 40 00
23 24 F4 FE 83 25 84 FE 03 25 C4 FE EF 00 00 18
93 07 05 00 23 22 F4 FE 83 27 44 FE 13 85 07 00
83 20 C1 01 03 24 81 01 13 01 01 02 67 80 00 00
13 01 01 FE 23 2E 11 00 23 2C 81 00 23 2A 91 00
13 04 01 02 B7 07 C0 00 93 87 47 00 83 A7 07 00
23 26 F4 FE 03 27 C4 FE 93 07 30 00 63 06 F7 0E
03 27 C4 FE 93 07 30 00 63 C4 E7 10 03 27 C4 FE
93 07 20 00 63 06 F7 0A 03 27 C4 FE 93 07 20 00
63 C8 E7 0E 83 27 C4 FE 63 8A 07 00 03 27 C4 FE
93 07 10 00 63 02 F7 06 6F 00 80 0D B7 17 40 00
93 84 07 F0 EF F0 DF E5 93 07 05 00 23 A0 F4 00
B7 07 C0 00 93 87 07 20 13 07 10 00 23 A0 E7 00
13 00 00 00 B7 07 C0 00 93 87 47 20 83 A7 07 00
E3 8A 07 FE B7 07 C0 00 93 87 87 20 83 A7 07 00
E3 82 07 FE B7 07 C0 00 93 87 C7 20 83 A7 07 00
E3 8A 07 FC 6F 00 C0 07 B7 17 40 00 93 84 47 F0
EF F0 DF E4 93 07 05 00 23 A0 F4 00 B7 07 C0 00
93 87 47 20 13 07 10 00 23 A0 E7 00 6F 00 00 00
B7 17 40 00 93 84 87 F0 EF F0 1F E7 93 07 05 00
23 A0 F4 00 B7 07 C0 00 93 87 87 20 13 07 10 00
23 A0 E7 00 6F 00 00 00 B7 17 40 00 93 84 C7 F0
EF F0 5F E9 93 07 05 00 23 A0 F4 00 B7 07 C0 00
93 87 C7 20 13 07 10 00 23 A0 E7 00 6F 00 00 00
13 00 00 00 13 85 07 00 83 20 C1 01 03 24 81 01
83 24 41 01 13 01 01 02 67 80 00 00 13 06 05 00
13 05 00 00 93 F6 15 00 63 84 06 00 33 05 C5 00
93 D5 15 00 13 16 16 00 E3 96 05 FE 67 80 00 00
