@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 13
@00000018
13 01 01 FB 23 26 81 04 13 04 01 05 93 07 10 00
23 2E F4 FA 93 07 50 00 23 20 F4 FC 93 07 70 00
23 22 F4 FC 93 07 30 00 23 24 F4 FC 93 07 50 00
23 26 F4 FC 93 07 90 00 23 28 F4 FC 93 07 20 03
23 2A F4 FC 93 07 20 00 23 2C F4 FC 93 07 90 00
23 20 F4 FE 23 26 04 FE 93 07 20 00 23 24 F4 FE
23 22 04 FE B7 17 40 00 93 87 07 F0 23 A0 07 00
6F 00 80 09 03 27 84 FE 83 27 C4 FE B3 07 F7 40
13 D7 F7 01 B3 07 F7 00 93 D7 17 40 13 87 07 00
83 27 C4 FE B3 87 E7 00 23 2E F4 FC 83 27 C4 FD
93 97 27 00 13 07 04 FF B3 07 F7 00 83 A7 C7 FC
03 27 04 FE 63 1E F7 00 93 07 10 00 23 22 F4 FE
B7 17 40 00 93 87 07 F0 13 07 10 00 23 A0 E7 00
83 27 C4 FD 93 97 27 00 13 07 04 FF B3 07 F7 00
83 A7 C7 FC 03 27 04 FE 63 DA E7 00 83 27 C4 FD
93 87 17 00 23 26 F4 FE 6F 00 00 01 83 27 C4 FD
93 87 F7 FF 23 24 F4 FE 03 27 C4 FE 83 27 84 FE
63 C6 E7 00 83 27 44 FE E3 8E 07 F4 13 00 00 00
13 85 07 00 03 24 C1 04 13 01 01 05 67 80 00 00
93 00 00 00 13 81 00 00 93 81 00 00 13 82 00 00
93 82 00 00 13 83 00 00 93 83 00 00 13 84 00 00
93 84 00 00 13 85 00 00 93 85 00 00 13 86 00 00
93 86 00 00 13 87 00 00 93 87 00 00 B7 02 C0 00
93 82 C2 00 03 A1 02 00 EF F0 9F E8
