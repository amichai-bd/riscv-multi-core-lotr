@00400800
02 00 00 00 03 00 00 00 04 00 00 00 0A 00 00 00
28 00 00 00
