@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 10 60 73 00 10 00
@000000A8
13 01 01 FD 23 26 81 02 13 04 01 03 23 2E A4 FC
23 2C B4 FC 23 2A C4 FC 03 27 84 FD 93 07 07 00
93 97 27 00 B3 87 E7 00 93 97 67 00 23 26 F4 FE
83 27 44 FD 93 97 27 00 23 24 F4 FE 03 27 84 FE
83 27 C4 FE 33 07 F7 00 B7 07 40 03 B3 07 F7 00
23 22 F4 FE 03 27 84 FE 83 27 C4 FE 33 07 F7 00
B7 07 40 03 93 87 07 14 B3 07 F7 00 23 20 F4 FE
83 27 C4 FD 13 97 27 00 B7 17 40 00 93 87 07 90
B3 07 F7 00 03 A7 07 00 83 27 44 FE 23 A0 E7 00
83 27 C4 FD 13 97 27 00 B7 17 40 00 93 87 07 A0
B3 07 F7 00 03 A7 07 00 83 27 04 FE 23 A0 E7 00
13 00 00 00 03 24 C1 02 13 01 01 03 67 80 00 00
13 01 01 FF 23 26 81 00 13 04 01 01 B7 17 40 00
93 87 07 98 23 A0 07 00 B7 17 40 00 93 87 07 A8
23 A0 07 00 B7 17 40 00 93 87 07 9C 37 47 62 52
13 07 07 C0 23 A0 E7 00 B7 17 40 00 93 87 07 AC
37 47 3C 00 13 07 A7 64 23 A0 E7 00 B7 17 40 00
93 87 47 9C 37 27 1C 1A 13 07 07 80 23 A0 E7 00
B7 17 40 00 93 87 47 AC 37 27 7E 00 13 07 87 81
23 A0 E7 00 B7 17 40 00 93 87 87 9C 37 47 42 40
13 07 07 C0 23 A0 E7 00 B7 17 40 00 93 87 87 AC
37 07 7E 00 13 07 C7 23 23 A0 E7 00 B7 17 40 00
93 87 C7 9C 37 47 42 40 13 07 07 C0 23 A0 E7 00
B7 17 40 00 93 87 C7 AC 37 47 3C 00 13 07 87 23
23 A0 E7 00 B7 17 40 00 93 87 07 9D 37 37 28 24
23 A0 E7 00 B7 17 40 00 93 87 07 AD 37 27 20 00
13 07 E7 07 23 A0 E7 00 B7 17 40 00 93 87 47 9D
37 87 02 3E 13 07 07 E0 23 A0 E7 00 B7 17 40 00
93 87 47 AD 37 47 3C 00 13 07 07 24 23 A0 E7 00
B7 17 40 00 93 87 87 9D 37 47 42 02 13 07 07 C0
23 A0 E7 00 B7 17 40 00 93 87 87 AD 37 47 3C 00
13 07 E7 23 23 A0 E7 00 B7 17 40 00 93 87 C7 9D
37 87 40 30 13 07 07 E0 23 A0 E7 00 B7 17 40 00
93 87 C7 AD 37 17 08 00 13 07 87 80 23 A0 E7 00
B7 17 40 00 93 87 07 9E 37 47 42 42 13 07 07 C0
23 A0 E7 00 B7 17 40 00 93 87 07 AE 37 47 3C 00
13 07 C7 23 23 A0 E7 00 B7 17 40 00 93 87 47 9E
37 47 42 42 13 07 07 C0 23 A0 E7 00 B7 17 40 00
93 87 47 AE 37 47 3E 00 13 07 C7 07 23 A0 E7 00
B7 17 40 00 93 87 47 A0 37 27 3C 66 13 07 07 80
23 A0 E7 00 B7 17 40 00 93 87 47 B0 37 87 66 00
13 07 67 E6 23 A0 E7 00 B7 17 40 00 93 87 C7 A0
37 47 3E 02 13 07 07 C0 23 A0 E7 00 B7 17 40 00
93 87 C7 B0 37 47 3C 00 13 07 27 E0 23 A0 E7 00
B7 17 40 00 93 87 47 A1 37 87 06 06 13 07 07 E0
23 A0 E7 00 B7 17 40 00 93 87 47 B1 37 07 7E 00
13 07 E7 67 23 A0 E7 00 B7 17 40 00 93 87 C7 A1
37 47 3E 02 13 07 07 C0 23 A0 E7 00 B7 17 40 00
93 87 C7 B1 37 27 3C 00 13 07 A7 23 23 A0 E7 00
B7 17 40 00 93 87 47 A3 37 47 66 5A 13 07 07 20
23 A0 E7 00 B7 17 40 00 93 87 47 B3 37 47 42 00
13 07 A7 25 23 A0 E7 00 B7 17 40 00 93 87 C7 A3
37 47 66 66 13 07 07 C0 23 A0 E7 00 B7 17 40 00
93 87 C7 B3 37 67 3C 00 13 07 67 66 23 A0 E7 00
B7 17 40 00 93 87 87 A4 37 47 66 66 13 07 07 E0
23 A0 E7 00 B7 17 40 00 93 87 87 B4 37 67 66 00
13 07 E7 63 23 A0 E7 00 B7 17 40 00 93 87 C7 A4
37 87 06 1E 13 07 07 C0 23 A0 E7 00 B7 17 40 00
93 87 C7 B4 37 67 3E 00 13 07 87 07 23 A0 E7 00
B7 17 40 00 93 87 07 A6 37 67 66 3C 13 07 07 60
23 A0 E7 00 B7 17 40 00 93 87 07 B6 37 67 66 00
13 07 C7 63 23 A0 E7 00 B7 17 40 00 93 87 C7 9A
13 07 F0 FF 23 A0 E7 00 B7 17 40 00 93 87 C7 AA
13 07 F0 FF 23 A0 E7 00 13 00 00 00 03 24 C1 00
13 01 01 01 67 80 00 00 13 01 01 FE 23 2E 11 00
23 2C 81 00 13 04 01 02 23 26 A4 FE 23 24 B4 FE
83 27 84 FE 93 87 67 00 13 86 07 00 83 25 C4 FE
13 05 70 04 EF F0 DF BC 83 27 84 FE 93 87 77 00
13 86 07 00 83 25 C4 FE 13 05 10 04 EF F0 5F BB
83 27 84 FE 93 87 87 00 13 86 07 00 83 25 C4 FE
13 05 D0 04 EF F0 DF B9 83 27 84 FE 93 87 97 00
13 86 07 00 83 25 C4 FE 13 05 50 04 EF F0 5F B8
83 27 84 FE 93 87 A7 00 13 86 07 00 83 25 C4 FE
13 05 00 02 EF F0 DF B6 83 27 84 FE 93 87 B7 00
13 86 07 00 83 25 C4 FE 13 05 30 05 EF F0 5F B5
83 27 84 FE 93 87 C7 00 13 86 07 00 83 25 C4 FE
13 05 30 04 EF F0 DF B3 83 27 84 FE 93 87 D7 00
13 86 07 00 83 25 C4 FE 13 05 F0 04 EF F0 5F B2
83 27 84 FE 93 87 E7 00 13 86 07 00 83 25 C4 FE
13 05 20 05 EF F0 DF B0 83 27 84 FE 93 87 F7 00
13 86 07 00 83 25 C4 FE 13 05 50 04 EF F0 5F AF
13 00 00 00 83 20 C1 01 03 24 81 01 13 01 01 02
67 80 00 00 13 01 01 FE 23 2E 11 00 23 2C 81 00
13 04 01 02 23 26 04 FE 6F 00 80 04 23 24 04 FE
6F 00 80 02 83 27 84 FE 93 97 17 00 03 26 C4 FE
93 85 07 00 13 05 00 02 EF F0 9F AA 83 27 84 FE
93 87 17 00 23 24 F4 FE 03 27 84 FE 93 07 B0 03
E3 DA E7 FC 83 27 C4 FE 93 87 17 00 23 26 F4 FE
03 27 C4 FE 93 07 F0 04 E3 DA E7 FA 13 00 00 00
13 00 00 00 83 20 C1 01 03 24 81 01 13 01 01 02
67 80 00 00 13 01 01 FE 23 2E 11 00 23 2C 81 00
13 04 01 02 23 26 04 FE 6F 00 00 03 03 26 C4 FE
93 05 00 00 13 05 B0 02 EF F0 9F A3 03 26 C4 FE
93 05 60 07 13 05 B0 02 EF F0 9F A2 83 27 C4 FE
93 87 17 00 23 26 F4 FE 03 27 C4 FE 93 07 F0 04
E3 D6 E7 FC 23 24 04 FE 6F 00 00 04 83 27 84 FE
93 97 17 00 13 06 00 00 93 85 07 00 13 05 B0 02
EF F0 1F 9F 83 27 84 FE 93 97 17 00 13 06 F0 04
93 85 07 00 13 05 B0 02 EF F0 9F 9D 83 27 84 FE
93 87 17 00 23 24 F4 FE 03 27 84 FE 93 07 B0 03
E3 DE E7 FA 13 00 00 00 13 00 00 00 83 20 C1 01
03 24 81 01 13 01 01 02 67 80 00 00 13 01 01 FE
23 2E 81 00 13 04 01 02 23 26 A4 FE 6F 00 00 01
83 27 C4 FE 93 87 F7 FF 23 26 F4 FE 83 27 C4 FE
E3 48 F0 FE 13 00 00 00 13 00 00 00 03 24 C1 01
13 01 01 02 67 80 00 00 13 01 01 FD 23 26 81 02
13 04 01 03 23 2E A4 FC B7 27 C0 03 93 87 C7 02
83 A7 07 00 23 26 F4 FE 03 27 C4 FE 93 07 10 00
63 08 F7 02 03 27 C4 FE 93 07 40 00 63 02 F7 02
03 27 C4 FE 93 07 80 00 63 0C F7 00 03 27 C4 FE
93 07 20 00 63 06 F7 00 83 27 C4 FD 23 26 F4 FE
03 27 C4 FD 93 07 10 00 63 1C F7 00 03 27 C4 FE
93 07 80 00 63 16 F7 00 83 27 C4 FD 23 26 F4 FE
03 27 C4 FD 93 07 80 00 63 1C F7 00 03 27 C4 FE
93 07 10 00 63 16 F7 00 83 27 C4 FD 23 26 F4 FE
03 27 C4 FD 93 07 40 00 63 1C F7 00 03 27 C4 FE
93 07 20 00 63 16 F7 00 83 27 C4 FD 23 26 F4 FE
03 27 C4 FD 93 07 20 00 63 1C F7 00 03 27 C4 FE
93 07 40 00 63 16 F7 00 83 27 C4 FD 23 26 F4 FE
83 27 C4 FE 13 85 07 00 03 24 C1 02 13 01 01 03
67 80 00 00 13 01 01 FD 23 26 81 02 13 04 01 03
23 2E A4 FC 23 2C B4 FC 23 2A C4 FC 23 28 D4 FC
83 27 04 FD 93 87 F7 FF 23 26 F4 FE 6F 00 80 07
03 27 C4 FE B7 07 00 40 93 87 F7 FF B3 07 F7 00
93 97 27 00 03 27 84 FD 33 07 F7 00 83 27 C4 FE
93 97 27 00 83 26 84 FD B3 87 F6 00 03 27 07 00
23 A0 E7 00 03 27 C4 FE B7 07 00 40 93 87 F7 FF
B3 07 F7 00 93 97 27 00 03 27 44 FD 33 07 F7 00
83 27 C4 FE 93 97 27 00 83 26 44 FD B3 87 F6 00
03 27 07 00 23 A0 E7 00 83 27 C4 FE 93 87 F7 FF
23 26 F4 FE 83 27 C4 FE E3 44 F0 F8 03 27 C4 FD
93 07 40 00 63 16 F7 02 83 27 84 FD 03 A7 47 00
83 27 84 FD 23 A0 E7 00 83 27 44 FD 93 87 47 00
83 A7 07 00 13 87 F7 FF 83 27 44 FD 23 A0 E7 00
03 27 C4 FD 93 07 20 00 63 16 F7 02 83 27 84 FD
03 A7 47 00 83 27 84 FD 23 A0 E7 00 83 27 44 FD
93 87 47 00 83 A7 07 00 13 87 17 00 83 27 44 FD
23 A0 E7 00 03 27 C4 FD 93 07 80 00 63 16 F7 02
83 27 84 FD 93 87 47 00 83 A7 07 00 13 87 F7 FF
83 27 84 FD 23 A0 E7 00 83 27 44 FD 03 A7 47 00
83 27 44 FD 23 A0 E7 00 03 27 C4 FD 93 07 10 00
63 16 F7 02 83 27 84 FD 93 87 47 00 83 A7 07 00
13 87 17 00 83 27 84 FD 23 A0 E7 00 83 27 44 FD
03 A7 47 00 83 27 44 FD 23 A0 E7 00 83 27 C4 FD
63 96 07 02 83 27 84 FD 93 87 47 00 83 A7 07 00
13 87 17 00 83 27 84 FD 23 A0 E7 00 83 27 44 FD
03 A7 47 00 83 27 44 FD 23 A0 E7 00 13 00 00 00
03 24 C1 02 13 01 01 03 67 80 00 00 13 01 01 FC
23 2E 11 02 23 2C 81 02 13 04 01 04 23 2E A4 FC
23 2C B4 FC 23 2A C4 FC 23 28 D4 FC 23 26 E4 FC
23 26 04 FE 6F 00 00 0F 83 27 C4 FE 93 97 27 00
03 27 84 FD B3 07 F7 00 83 A7 07 00 63 86 07 0C
83 27 C4 FE 93 97 27 00 03 27 04 FD B3 07 F7 00
83 A7 07 00 93 96 17 00 83 27 C4 FE 93 97 27 00
03 27 44 FD B3 07 F7 00 83 A7 07 00 13 86 07 00
93 85 06 00 13 05 B0 02 EF F0 8F E4 83 27 C4 FE
93 87 17 00 93 97 27 00 03 27 84 FD B3 07 F7 00
83 A7 07 00 63 9A 07 06 83 27 C4 FD 63 84 07 02
83 27 C4 FE 93 87 17 00 93 97 27 00 03 27 84 FD
B3 07 F7 00 13 07 10 00 23 A0 E7 00 23 2E 04 FC
6F 00 80 04 83 27 C4 FE 93 87 17 00 93 97 27 00
03 27 04 FD B3 07 F7 00 83 A7 07 00 93 96 17 00
83 27 C4 FE 93 87 17 00 93 97 27 00 03 27 44 FD
B3 07 F7 00 83 A7 07 00 13 86 07 00 93 85 06 00
13 05 00 02 EF F0 CF DB 83 27 C4 FE 93 87 17 00
23 26 F4 FE 03 27 C4 FE 83 27 C4 FC E3 46 F7 F0
13 00 00 00 13 00 00 00 83 20 C1 03 03 24 81 03
13 01 01 04 67 80 00 00 13 01 01 FC 23 2E 81 02
13 04 01 04 23 2E A4 FC 23 2C B4 FC 23 2A C4 FC
23 28 D4 FC 23 26 E4 FC 23 24 F4 FC 03 27 84 FD
83 27 04 FD 63 1C F7 00 03 27 44 FD 83 27 C4 FC
63 16 F7 00 93 07 10 00 6F 00 80 00 93 07 00 00
23 26 F4 FE 83 27 C4 FE 63 8C 07 00 83 27 84 FC
83 A7 07 00 13 87 17 00 83 27 84 FC 23 A0 E7 00
83 27 C4 FE 13 85 07 00 03 24 C1 03 13 01 01 04
67 80 00 00 13 01 01 FD 23 26 81 02 13 04 01 03
23 2E A4 FC 23 2C B4 FC 23 26 04 FE 83 27 C4 FD
63 96 07 00 93 07 10 00 23 26 F4 FE 03 27 C4 FD
93 07 F0 04 63 16 F7 00 93 07 10 00 23 26 F4 FE
83 27 84 FD 63 96 07 00 93 07 10 00 23 26 F4 FE
03 27 84 FD 93 07 B0 03 63 16 F7 00 93 07 10 00
23 26 F4 FE 83 27 C4 FE 13 85 07 00 03 24 C1 02
13 01 01 03 67 80 00 00 13 01 01 FE 23 2E 11 00
23 2C 81 00 13 04 01 02 23 26 A4 FE 23 24 B4 FE
83 27 84 FE 83 A7 07 00 93 05 30 00 13 85 07 00
EF 00 40 2C 93 07 05 00 13 87 07 00 83 27 C4 FE
83 A7 07 00 93 85 07 00 13 05 07 00 EF 00 40 28
93 07 05 00 13 87 07 00 93 57 F7 41 93 D7 A7 01
33 07 F7 00 13 77 F7 03 B3 07 F7 40 13 87 17 00
83 27 C4 FE 23 A0 E7 00 83 27 C4 FE 83 A7 07 00
13 D7 F7 41 13 77 37 00 B3 07 F7 00 93 D7 27 40
13 87 07 00 83 27 84 FE 83 A7 07 00 93 85 07 00
13 05 07 00 EF 00 C0 22 93 07 05 00 13 87 07 00
93 57 F7 41 93 D7 B7 01 33 07 F7 00 13 77 F7 01
B3 07 F7 40 13 87 17 00 83 27 84 FE 23 A0 E7 00
13 00 00 00 83 20 C1 01 03 24 81 01 13 01 01 02
67 80 00 00 13 01 01 F1 23 26 11 0E 23 24 81 0E
13 04 01 0F 93 07 10 00 23 26 F4 FE 93 07 50 00
23 22 F4 F2 93 07 50 00 23 20 F4 F2 23 2E 04 F0
23 24 04 FE 23 22 04 FE EF F0 DF 92 23 20 04 FE
6F 00 80 06 83 27 04 FE 13 87 47 01 83 27 04 FE
93 97 27 00 93 87 07 FF B3 87 87 00 23 A8 E7 FA
83 27 04 FE 93 97 27 00 93 87 07 FF B3 87 87 00
13 07 40 01 23 AA E7 F6 83 27 04 FE 93 A7 57 00
93 F7 F7 0F 13 87 07 00 83 27 04 FE 93 97 27 00
93 87 07 FF B3 87 87 00 23 AC E7 F2 83 27 04 FE
93 87 17 00 23 20 F4 FE 03 27 04 FE 93 07 E0 00
E3 DA E7 F8 03 25 C4 FE EF F0 1F 9A 23 26 A4 FE
83 27 44 FE 63 90 07 02 13 07 44 F6 93 07 04 FA
93 06 F0 00 13 06 07 00 93 85 07 00 03 25 C4 FE
EF F0 5F A6 83 25 04 FA 03 26 44 F6 83 26 44 F2
03 27 04 F2 93 07 C4 F1 13 05 84 F2 EF F0 DF D3
23 2E A4 FC 03 27 C4 FD 93 07 10 00 63 12 F7 02
13 07 04 F2 93 07 44 F2 93 05 07 00 13 85 07 00
EF F0 9F E0 83 27 84 FE 93 87 17 00 23 24 F4 FE
93 05 40 01 13 05 30 00 EF F0 0F E9 83 27 04 F2
93 97 17 00 03 27 44 F2 13 06 07 00 93 85 07 00
13 05 F0 04 EF F0 CF A6 93 06 44 F6 13 06 04 FA
93 07 84 F2 13 07 F0 00 93 85 07 00 03 25 C4 FD
EF F0 DF B8 83 27 84 FE 93 87 07 03 13 06 70 02
93 05 30 00 13 85 07 00 EF F0 8F A3 83 27 04 FA
03 27 44 F6 93 05 07 00 13 85 07 00 EF F0 9F D1
23 22 A4 FE 23 2E 04 FC B7 57 00 00 13 85 07 E2
EF F0 DF 86 6F F0 1F F0 13 01 01 FE 23 2E 11 00
23 2C 81 00 13 04 01 02 B7 07 C0 00 83 A7 07 00
23 26 F4 FE EF F0 CF AA EF F0 CF F0 03 27 C4 FE
93 07 40 00 63 14 F7 00 EF F0 DF E1 6F 00 00 00
13 06 05 00 13 05 00 00 93 F6 15 00 63 84 06 00
33 05 C5 00 93 D5 15 00 13 16 16 00 E3 96 05 FE
67 80 00 00 63 40 05 06 63 C6 05 06 13 86 05 00
93 05 05 00 13 05 F0 FF 63 0C 06 02 93 06 10 00
63 7A B6 00 63 58 C0 00 13 16 16 00 93 96 16 00
E3 6A B6 FE 13 05 00 00 63 E6 C5 00 B3 85 C5 40
33 65 D5 00 93 D6 16 00 13 56 16 00 E3 96 06 FE
67 80 00 00 93 82 00 00 EF F0 5F FB 13 85 05 00
67 80 02 00 33 05 A0 40 63 48 B0 00 B3 05 B0 40
6F F0 DF F9 B3 05 B0 40 93 82 00 00 EF F0 1F F9
33 05 A0 40 67 80 02 00 93 82 00 00 63 CA 05 00
63 4C 05 00 EF F0 9F F7 13 85 05 00 67 80 02 00
B3 05 B0 40 E3 58 05 FE 33 05 A0 40 EF F0 1F F6
33 05 B0 40 67 80 02 00
