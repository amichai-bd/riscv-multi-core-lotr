@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 80 04 67 80 00 00
@0000001C
13 01 01 FE 23 2E 81 00 13 04 01 02 93 07 50 00
23 26 F4 FE 93 07 40 00 23 24 F4 FE 03 27 C4 FE
83 27 84 FE B3 07 F7 00 23 22 F4 FE 13 00 00 00
13 85 07 00 03 24 C1 01 13 01 01 02 67 80 00 00
93 00 00 00 13 81 00 00 93 81 00 00 13 82 00 00
93 82 00 00 13 83 00 00 93 83 00 00 13 84 00 00
93 84 00 00 13 85 00 00 93 85 00 00 13 86 00 00
93 86 00 00 13 87 00 00 93 87 00 00 B7 02 C0 00
93 82 C2 00 03 A1 02 00 EF F0 9F F7
