@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 C0 0C 73 00 10 00
@000000A8
13 01 01 FD 23 26 81 02 13 04 01 03 23 2E A4 FC
23 2C B4 FC 23 2A C4 FC 23 28 D4 FC 6F 00 80 08
03 27 44 FD 83 27 84 FD B3 07 F7 40 13 D7 F7 01
B3 07 F7 00 93 D7 17 40 13 87 07 00 83 27 84 FD
B3 87 E7 00 23 26 F4 FE 83 27 C4 FE 93 97 27 00
03 27 C4 FD B3 07 F7 00 83 A7 07 00 03 27 04 FD
63 16 F7 00 83 27 C4 FE 6F 00 C0 04 83 27 C4 FE
93 97 27 00 03 27 C4 FD B3 07 F7 00 83 A7 07 00
03 27 04 FD 63 DA E7 00 83 27 C4 FE 93 87 17 00
23 2C F4 FC 6F 00 00 01 83 27 C4 FE 93 87 F7 FF
23 2A F4 FC 03 27 84 FD 83 27 44 FD E3 DA E7 F6
93 07 F0 FF 13 85 07 00 03 24 C1 02 13 01 01 03
67 80 00 00 13 01 01 FD 23 26 11 02 23 24 81 02
13 04 01 03 B7 17 40 00 93 87 07 80 83 A5 07 00
03 A6 47 00 83 A6 87 00 03 A7 C7 00 83 A7 07 01
23 28 B4 FC 23 2A C4 FC 23 2C D4 FC 23 2E E4 FC
23 20 F4 FE 93 07 60 00 23 26 F4 FE 93 07 A0 00
23 24 F4 FE 83 27 C4 FE 13 87 F7 FF 93 07 04 FD
83 26 84 FE 13 06 07 00 93 05 00 00 13 85 07 00
EF F0 1F ED 23 22 A4 FE 03 27 44 FE 93 07 F0 FF
63 1A F7 00 B7 17 40 00 93 87 07 F0 23 A0 07 00
6F 00 40 01 B7 17 40 00 93 87 07 F0 13 07 10 00
23 A0 E7 00 93 07 00 00 13 85 07 00 83 20 C1 02
03 24 81 02 13 01 01 03 67 80 00 00
