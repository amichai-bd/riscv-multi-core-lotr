@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 80 26 73 00 10 00
@000000A8
13 01 01 FD 23 26 81 02 13 04 01 03 23 2E A4 FC
23 2C B4 FC 83 27 C4 FD 83 A7 07 00 23 26 F4 FE
83 27 84 FD 03 A7 07 00 83 27 C4 FD 23 A0 E7 00
03 27 C4 FE 83 27 84 FD 23 A0 E7 00 13 00 00 00
03 24 C1 02 13 01 01 03 67 80 00 00 13 01 01 FD
23 26 11 02 23 24 81 02 13 04 01 03 23 2E A4 FC
23 2C B4 FC 23 26 04 FE 6F 00 C0 09 23 24 04 FE
6F 00 00 07 83 27 84 FE 93 97 27 00 03 27 C4 FD
B3 07 F7 00 03 A7 07 00 83 27 84 FE 93 87 17 00
93 97 27 00 83 26 C4 FD B3 87 F6 00 83 A7 07 00
63 DA E7 02 83 27 84 FE 93 97 27 00 03 27 C4 FD
B3 06 F7 00 83 27 84 FE 93 87 17 00 93 97 27 00
03 27 C4 FD B3 07 F7 00 93 85 07 00 13 85 06 00
EF F0 1F F3 83 27 84 FE 93 87 17 00 23 24 F4 FE
03 27 84 FD 83 27 C4 FE B3 07 F7 40 93 87 F7 FF
03 27 84 FE E3 40 F7 F8 83 27 C4 FE 93 87 17 00
23 26 F4 FE 83 27 84 FD 93 87 F7 FF 03 27 C4 FE
E3 4E F7 F4 13 00 00 00 13 00 00 00 83 20 C1 02
03 24 81 02 13 01 01 03 67 80 00 00 13 01 01 FC
23 2E 81 02 13 04 01 04 23 26 A4 FC 23 24 B4 FC
23 22 C4 FC 83 27 44 FC 13 07 F0 0F 23 A0 E7 00
83 27 44 FC 93 87 47 00 13 07 E0 0F 23 A0 E7 00
23 26 04 FE 6F 00 C0 0D 23 24 04 FE 6F 00 C0 0B
83 27 44 FC 93 87 C7 00 13 07 E0 0F 23 A0 E7 00
23 2E 04 FC 23 22 04 FE 6F 00 C0 04 83 27 C4 FE
13 97 27 00 83 27 44 FE B3 07 F7 00 93 97 27 00
03 27 C4 FC B3 07 F7 00 83 A7 07 00 23 20 F4 FE
83 27 44 FC 93 87 87 01 83 26 04 FE 03 27 84 FD
33 87 E6 00 23 A0 E7 00 83 27 44 FE 93 87 17 00
23 22 F4 FE 03 27 44 FE 93 07 30 00 E3 D8 E7 FA
83 27 44 FC 93 87 C7 01 83 26 04 FE 03 27 84 FD
33 87 E6 00 23 A0 E7 00 83 27 C4 FE 13 97 27 00
83 27 84 FE B3 07 F7 00 93 97 27 00 03 27 44 FC
B3 07 F7 00 03 27 C4 FD 23 A0 E7 00 83 27 84 FE
93 87 17 00 23 24 F4 FE 03 27 84 FE 93 07 30 00
E3 D0 E7 F4 83 27 C4 FE 93 87 17 00 23 26 F4 FE
03 27 C4 FE 93 07 30 00 E3 D0 E7 F2 13 00 00 00
13 00 00 00 03 24 C1 03 13 01 01 04 67 80 00 00
13 01 01 F4 23 2E 11 0A 23 2C 81 0A 13 04 01 0C
B7 07 C0 00 83 A7 07 00 23 20 F4 FE 23 2E 04 FC
83 27 04 FE 93 87 C7 FF 13 07 70 00 63 60 F7 2E
13 97 27 00 B7 17 40 00 93 87 07 8C B3 07 F7 00
83 A7 07 00 67 80 07 00 B7 07 C0 01 93 87 07 15
23 A0 07 00 B7 17 40 02 93 87 07 90 23 22 F4 FC
93 05 80 00 03 25 44 FC EF F0 5F D8 6F 00 00 00
B7 17 40 00 93 87 07 80 83 A8 07 00 03 A8 47 00
03 A5 87 00 83 A5 C7 00 03 A6 07 01 83 A6 47 01
03 A7 87 01 83 A7 C7 01 23 22 14 F9 23 24 04 F9
23 26 A4 F8 23 28 B4 F8 23 2A C4 F8 23 2C D4 F8
23 2E E4 F8 23 20 F4 FA 23 26 04 FE 6F 00 C0 03
83 27 C4 FE 13 97 27 00 B7 17 40 00 93 87 07 90
33 07 F7 00 83 27 C4 FE 93 97 27 00 93 06 04 FF
B3 87 F6 00 83 A7 47 F9 23 20 F7 00 83 27 C4 FE
93 87 17 00 23 26 F4 FE 03 27 C4 FE 93 07 70 00
E3 D0 E7 FC B7 07 C0 02 93 87 47 15 13 07 10 00
23 A0 E7 00 6F 00 00 00 23 24 04 FC B7 17 40 00
13 87 07 82 93 07 44 F4 93 06 07 00 13 07 00 04
13 06 07 00 93 85 06 00 13 85 07 00 EF 00 80 1E
B7 17 40 00 13 87 07 86 93 07 44 F8 93 06 07 00
13 07 00 04 13 06 07 00 93 85 06 00 13 85 07 00
EF 00 40 1C 23 24 04 FE 6F 00 80 06 83 27 84 FE
13 97 27 00 B7 17 40 00 93 87 07 A0 33 07 F7 00
83 27 84 FE 93 97 27 00 93 06 04 FF B3 87 F6 00
83 A7 47 F5 23 20 F7 00 83 27 84 FE 13 97 27 00
B7 17 40 00 93 87 07 B0 33 07 F7 00 83 27 84 FE
93 97 27 00 93 06 04 FF B3 87 F6 00 83 A7 47 F9
23 20 F7 00 83 27 84 FE 93 87 17 00 23 24 F4 FE
03 27 84 FE 93 07 F0 00 E3 DA E7 F8 B7 07 C0 02
93 87 87 15 13 07 10 00 23 A0 E7 00 6F 00 00 00
6F 00 00 00 B7 17 40 00 93 87 07 8A 83 A8 07 00
03 A8 47 00 03 A5 87 00 83 A5 C7 00 03 A6 07 01
83 A6 47 01 03 A7 87 01 83 A7 C7 01 23 22 14 F9
23 24 04 F9 23 26 A4 F8 23 28 B4 F8 23 2A C4 F8
23 2C D4 F8 23 2E E4 F8 23 20 F4 FA 23 22 04 FE
6F 00 C0 03 83 27 44 FE 13 97 27 00 B7 17 40 00
93 87 07 90 33 07 F7 00 83 27 44 FE 93 97 27 00
93 06 04 FF B3 87 F6 00 83 A7 47 F9 23 20 F7 00
83 27 44 FE 93 87 17 00 23 22 F4 FE 03 27 44 FE
93 07 70 00 E3 D0 E7 FC B7 07 C0 01 93 87 07 15
13 07 10 00 23 A0 E7 00 6F 00 00 00 B7 07 C0 02
93 87 47 15 23 A0 07 00 B7 17 40 01 93 87 07 90
23 26 F4 FC 93 05 80 00 03 25 C4 FC EF F0 1F B3
6F 00 00 00 B7 07 C0 02 93 87 87 15 23 A0 07 00
B7 17 40 01 93 87 07 A0 23 2C F4 FC B7 17 40 01
93 87 07 B0 23 2A F4 FC B7 17 40 01 93 87 07 C0
23 28 F4 FC 03 26 04 FD 83 25 44 FD 03 25 84 FD
EF F0 DF BC 6F 00 80 00 6F 00 00 00 93 07 00 00
13 85 07 00 83 20 C1 0B 03 24 81 0B 13 01 01 0C
67 80 00 00 B3 C7 A5 00 93 F7 37 00 B3 08 C5 00
63 96 07 06 93 07 30 00 63 F2 C7 06 93 77 35 00
13 07 05 00 63 9A 07 0C 13 F6 C8 FF B3 06 E6 40
93 07 00 02 93 02 00 02 63 C2 D7 06 93 86 05 00
93 07 07 00 63 78 C7 02 03 A8 06 00 93 87 47 00
93 86 46 00 23 AE 07 FF E3 E8 C7 FE 93 07 F6 FF
B3 87 E7 40 93 F7 C7 FF 93 87 47 00 33 07 F7 00
B3 85 F5 00 63 68 17 01 67 80 00 00 13 07 05 00
E3 7C 15 FF 83 C7 05 00 13 07 17 00 93 85 15 00
A3 0F F7 FE E3 68 17 FF 67 80 00 00 83 A6 45 00
83 A7 C5 01 83 AF 05 00 03 AF 85 00 83 AE C5 00
03 AE 05 01 03 A3 45 01 03 A8 85 01 23 22 D7 00
83 A6 05 02 23 20 F7 01 23 24 E7 01 23 26 D7 01
23 28 C7 01 23 2A 67 00 23 2C 07 01 23 2E F7 00
13 07 47 02 B3 07 E6 40 23 2E D7 FE 93 85 45 02
E3 C6 F2 FA 6F F0 9F F4 83 C6 05 00 13 07 17 00
93 77 37 00 A3 0F D7 FE 93 85 15 00 E3 8E 07 F0
83 C6 05 00 13 07 17 00 93 77 37 00 A3 0F D7 FE
93 85 15 00 E3 9A 07 FC 6F F0 1F F0
@00400800
0C 00 00 00 02 00 00 00 00 00 00 00 06 00 00 00
0A 00 00 00 12 00 00 00 64 00 00 00 04 00 00 00
01 00 00 00 02 00 00 00 03 00 00 00 04 00 00 00
05 00 00 00 06 00 00 00 07 00 00 00 08 00 00 00
09 00 00 00 0A 00 00 00 0B 00 00 00 0C 00 00 00
14 00 00 00 0E 00 00 00 0F 00 00 00 10 00 00 00
0D 00 00 00 0E 00 00 00 0F 00 00 00 10 00 00 00
09 00 00 00 0A 00 00 00 0B 00 00 00 0C 00 00 00
05 00 00 00 06 00 00 00 07 00 00 00 08 00 00 00
01 00 00 00 02 00 00 00 03 00 00 00 04 00 00 00
06 00 00 00 01 00 00 00 00 00 00 00 03 00 00 00
05 00 00 00 09 00 00 00 32 00 00 00 02 00 00 00
50 03 00 00 78 03 00 00 20 04 00 00 F8 04 00 00
FC 04 00 00 A4 05 00 00 CC 05 00 00 10 06 00 00
