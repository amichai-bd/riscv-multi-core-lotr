//-----------------------------------------------------------------------------
// Title            : Lotar 
// Project          : LOTR: Lord-Of-The-Ring
//-----------------------------------------------------------------------------
// File             : lotr.sv 
// Original Author  : Amichai
// Created          : 5/2021
//-----------------------------------------------------------------------------
// Description :
// 
//
// 
//------------------------------------------------------------------------------
// Modification history :
//
//
//------------------------------------------------------------------------------

`include "lotr_defines.sv"
module lotr
    import lotr_pkg::*;  
    (
    //General Interface
    input   logic        QClk                   ,
    input   logic        RstQnnnH               ,
    );

//=========================================
//=====    ===========
//=========================================



endmodule // module lotr
