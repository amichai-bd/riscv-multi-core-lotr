@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 90 34 73 00 10 00
@000000A8
13 01 01 FD 23 26 81 02 13 04 01 03 23 2E A4 FC
23 2C B4 FC 23 2A C4 FC 03 27 84 FD 93 07 07 00
93 97 27 00 B3 87 E7 00 93 97 67 00 23 26 F4 FE
83 27 44 FD 93 97 27 00 23 24 F4 FE 03 27 84 FE
83 27 C4 FE 33 07 F7 00 B7 07 40 03 B3 07 F7 00
23 22 F4 FE 03 27 84 FE 83 27 C4 FE 33 07 F7 00
B7 07 40 03 93 87 07 14 B3 07 F7 00 23 20 F4 FE
83 27 C4 FD 13 97 27 00 B7 17 40 00 93 87 07 90
B3 07 F7 00 03 A7 07 00 83 27 44 FE 23 A0 E7 00
83 27 C4 FD 13 97 27 00 B7 17 40 00 93 87 07 A0
B3 07 F7 00 03 A7 07 00 83 27 04 FE 23 A0 E7 00
13 00 00 00 03 24 C1 02 13 01 01 03 67 80 00 00
13 01 01 FD 23 26 11 02 23 24 81 02 13 04 01 03
23 2E A4 FC 23 26 04 FE 23 24 04 FE 23 22 04 FE
B7 07 C0 00 93 87 07 20 83 A7 07 00 23 22 F4 FE
B7 07 C0 00 93 87 47 20 83 A7 07 00 23 24 F4 FE
6F 00 00 0C 83 27 C4 FE 93 97 27 00 03 27 C4 FD
B3 07 F7 00 03 A7 07 00 93 07 A0 00 63 1A F7 02
23 22 04 FE 83 27 84 FE 93 87 27 00 23 24 F4 FE
03 27 84 FE 93 07 80 07 63 14 F7 00 23 24 04 FE
83 27 C4 FE 93 87 17 00 23 26 F4 FE 6F 00 40 07
83 27 C4 FE 93 97 27 00 03 27 C4 FD B3 07 F7 00
83 A7 07 00 03 27 84 FE 83 26 44 FE 13 86 06 00
93 05 07 00 13 85 07 00 EF F0 9F E8 83 27 44 FE
93 87 17 00 23 22 F4 FE 03 27 44 FE 93 07 00 05
63 12 F7 02 23 22 04 FE 83 27 84 FE 93 87 27 00
23 24 F4 FE 03 27 84 FE 93 07 80 07 63 14 F7 00
23 24 04 FE 83 27 C4 FE 93 87 17 00 23 26 F4 FE
83 27 C4 FE 93 97 27 00 03 27 C4 FD B3 07 F7 00
83 A7 07 00 E3 98 07 F2 B7 07 C0 00 93 87 07 20
03 27 44 FE 23 A0 E7 00 B7 07 C0 00 93 87 47 20
03 27 84 FE 23 A0 E7 00 13 00 00 00 83 20 C1 02
03 24 81 02 13 01 01 03 67 80 00 00 13 01 01 FF
23 26 81 00 13 04 01 01 B7 17 40 00 93 87 47 A0
37 27 3C 66 13 07 07 80 23 A0 E7 00 B7 17 40 00
93 87 47 B0 37 87 66 00 13 07 67 E6 23 A0 E7 00
B7 17 40 00 93 87 87 A0 37 27 22 3E 13 07 07 E0
23 A0 E7 00 B7 17 40 00 93 87 87 B0 37 27 1E 00
13 07 E7 23 23 A0 E7 00 B7 17 40 00 93 87 07 98
23 A0 07 00 B7 17 40 00 93 87 07 A8 23 A0 07 00
B7 17 40 00 93 87 07 9B 23 A0 07 00 B7 17 40 00
93 87 07 AB 37 27 1E 06 13 07 87 81 23 A0 E7 00
B7 17 40 00 93 87 87 9B 23 A0 07 00 B7 17 40 00
93 87 87 AB 37 27 18 00 13 07 07 80 23 A0 E7 00
B7 17 40 00 93 87 07 9C 37 47 62 52 13 07 07 C0
23 A0 E7 00 B7 17 40 00 93 87 07 AC 37 47 3C 00
13 07 A7 64 23 A0 E7 00 B7 17 40 00 93 87 47 9C
37 27 1C 1A 13 07 07 80 23 A0 E7 00 B7 17 40 00
93 87 47 AC 37 27 7E 00 13 07 87 81 23 A0 E7 00
B7 17 40 00 93 87 87 9C 37 47 42 40 13 07 07 C0
23 A0 E7 00 B7 17 40 00 93 87 87 AC 37 07 7E 00
13 07 C7 23 23 A0 E7 00 B7 17 40 00 93 87 C7 9C
37 47 42 40 13 07 07 C0 23 A0 E7 00 B7 17 40 00
93 87 C7 AC 37 47 3C 00 13 07 87 23 23 A0 E7 00
B7 17 40 00 93 87 07 9D 37 37 28 24 23 A0 E7 00
B7 17 40 00 93 87 07 AD 37 27 20 00 13 07 E7 07
23 A0 E7 00 B7 17 40 00 93 87 47 9D 37 87 02 3E
13 07 07 E0 23 A0 E7 00 B7 17 40 00 93 87 47 AD
37 47 3C 00 13 07 07 24 23 A0 E7 00 B7 17 40 00
93 87 87 9D 37 47 42 02 13 07 07 C0 23 A0 E7 00
B7 17 40 00 93 87 87 AD 37 47 3C 00 13 07 E7 23
23 A0 E7 00 B7 17 40 00 93 87 C7 9D 37 87 40 30
13 07 07 E0 23 A0 E7 00 B7 17 40 00 93 87 C7 AD
37 17 08 00 13 07 87 80 23 A0 E7 00 B7 17 40 00
93 87 07 9E 37 47 42 42 13 07 07 C0 23 A0 E7 00
B7 17 40 00 93 87 07 AE 37 47 3C 00 13 07 C7 23
23 A0 E7 00 B7 17 40 00 93 87 47 9E 37 47 42 42
13 07 07 C0 23 A0 E7 00 B7 17 40 00 93 87 47 AE
37 47 3E 00 13 07 C7 07 23 A0 E7 00 B7 17 40 00
93 87 47 A0 37 27 3C 66 13 07 07 80 23 A0 E7 00
B7 17 40 00 93 87 47 B0 37 87 66 00 13 07 67 E6
23 A0 E7 00 B7 17 40 00 93 87 87 A0 37 27 22 3E
13 07 07 E0 23 A0 E7 00 B7 17 40 00 93 87 87 B0
37 27 1E 00 13 07 E7 23 23 A0 E7 00 B7 17 40 00
93 87 C7 A0 37 47 3E 02 13 07 07 C0 23 A0 E7 00
B7 17 40 00 93 87 C7 B0 37 47 3C 00 13 07 27 E0
23 A0 E7 00 B7 17 40 00 93 87 07 A1 37 27 3E 22
13 07 07 E0 23 A0 E7 00 B7 17 40 00 93 87 07 B1
37 47 1E 00 13 07 27 E2 23 A0 E7 00 B7 17 40 00
93 87 47 A1 37 87 06 06 13 07 07 E0 23 A0 E7 00
B7 17 40 00 93 87 47 B1 37 07 7E 00 13 07 E7 67
23 A0 E7 00 B7 17 40 00 93 87 87 A1 37 87 06 06
13 07 07 E0 23 A0 E7 00 B7 17 40 00 93 87 87 B1
37 07 06 00 13 07 E7 67 23 A0 E7 00 B7 17 40 00
93 87 C7 A1 37 47 3E 02 13 07 07 C0 23 A0 E7 00
B7 17 40 00 93 87 C7 B1 37 27 3C 00 13 07 A7 23
23 A0 E7 00 B7 17 40 00 93 87 07 A2 37 67 66 66
13 07 07 60 23 A0 E7 00 B7 17 40 00 93 87 07 B2
37 67 66 00 13 07 E7 67 23 A0 E7 00 B7 17 40 00
93 87 47 A2 37 87 18 18 13 07 07 E0 23 A0 E7 00
B7 17 40 00 93 87 47 B2 37 27 7E 00 13 07 87 81
23 A0 E7 00 B7 17 40 00 93 87 87 A2 37 67 60 60
23 A0 E7 00 B7 17 40 00 93 87 87 B2 37 67 7C 00
13 07 67 66 23 A0 E7 00 B7 17 40 00 93 87 C7 A2
37 47 66 3E 13 07 07 60 23 A0 E7 00 B7 17 40 00
93 87 C7 B2 37 67 46 00 13 07 E7 63 23 A0 E7 00
B7 17 40 00 93 87 07 A3 37 07 06 06 13 07 07 60
23 A0 E7 00 B7 17 40 00 93 87 07 B3 37 07 7E 00
13 07 67 60 23 A0 E7 00 B7 17 40 00 93 87 47 A3
37 47 66 5A 13 07 07 20 23 A0 E7 00 B7 17 40 00
93 87 47 B3 37 47 42 00 13 07 A7 25 23 A0 E7 00
B7 17 40 00 93 87 87 A3 37 67 66 6E 13 07 07 20
23 A0 E7 00 B7 17 40 00 93 87 87 B3 37 67 46 00
13 07 67 67 23 A0 E7 00 B7 17 40 00 93 87 C7 A3
37 47 66 66 13 07 07 C0 23 A0 E7 00 B7 17 40 00
93 87 C7 B3 37 67 3C 00 13 07 67 66 23 A0 E7 00
B7 17 40 00 93 87 07 A4 37 47 66 66 13 07 07 E0
23 A0 E7 00 B7 17 40 00 93 87 07 B4 37 07 06 00
13 07 E7 63 23 A0 E7 00 B7 17 40 00 93 87 47 A4
37 47 42 42 13 07 07 C0 23 A0 E7 00 B7 17 40 00
93 87 47 B4 37 67 7C 00 13 07 27 25 23 A0 E7 00
B7 17 40 00 93 87 87 A4 37 47 66 66 13 07 07 E0
23 A0 E7 00 B7 17 40 00 93 87 87 B4 37 67 66 00
13 07 E7 63 23 A0 E7 00 B7 17 40 00 93 87 C7 A4
37 87 06 1E 13 07 07 C0 23 A0 E7 00 B7 17 40 00
93 87 C7 B4 37 67 3E 00 13 07 87 07 23 A0 E7 00
B7 17 40 00 93 87 07 A5 37 87 18 18 13 07 07 E0
23 A0 E7 00 B7 17 40 00 93 87 07 B5 37 27 18 00
13 07 87 81 23 A0 E7 00 B7 17 40 00 93 87 47 A5
37 67 66 66 13 07 07 60 23 A0 E7 00 B7 17 40 00
93 87 47 B5 37 87 3C 00 13 07 67 E6 23 A0 E7 00
B7 17 40 00 93 87 87 A5 37 67 66 66 13 07 07 60
23 A0 E7 00 B7 17 40 00 93 87 87 B5 37 47 18 00
13 07 67 C6 23 A0 E7 00 B7 17 40 00 93 87 C7 A5
37 47 42 42 13 07 07 20 23 A0 E7 00 B7 17 40 00
93 87 C7 B5 37 87 42 00 13 07 A7 E5 23 A0 E7 00
B7 17 40 00 93 87 07 A6 37 67 66 3C 13 07 07 60
23 A0 E7 00 B7 17 40 00 93 87 07 B6 37 67 66 00
13 07 C7 63 23 A0 E7 00 B7 17 40 00 93 87 47 A6
37 67 66 3C 13 07 07 60 23 A0 E7 00 B7 17 40 00
93 87 47 B6 37 27 18 00 13 07 87 81 23 A0 E7 00
B7 17 40 00 93 87 87 A6 37 87 20 10 13 07 07 E0
23 A0 E7 00 B7 17 40 00 93 87 87 B6 37 07 7E 00
13 07 87 40 23 A0 E7 00 B7 17 40 00 93 87 C7 AA
13 07 F0 FF 23 A0 E7 00 13 00 00 00 03 24 C1 00
13 01 01 01 67 80 00 00 13 01 01 FE 23 2E 11 00
23 2C 81 00 13 04 01 02 23 26 A4 FE 13 06 50 00
83 25 C4 FE 13 05 80 04 EF F0 8F F6 13 06 60 00
83 25 C4 FE 13 05 50 04 EF F0 8F F5 13 06 70 00
83 25 C4 FE 13 05 C0 04 EF F0 8F F4 13 06 80 00
83 25 C4 FE 13 05 C0 04 EF F0 8F F3 13 06 90 00
83 25 C4 FE 13 05 F0 04 EF F0 8F F2 13 06 A0 00
83 25 C4 FE 13 05 00 02 EF F0 8F F1 13 06 B0 00
83 25 C4 FE 13 05 70 05 EF F0 8F F0 13 06 C0 00
83 25 C4 FE 13 05 F0 04 EF F0 8F EF 13 06 D0 00
83 25 C4 FE 13 05 20 05 EF F0 8F EE 13 06 E0 00
83 25 C4 FE 13 05 C0 04 EF F0 8F ED 13 06 F0 00
83 25 C4 FE 13 05 40 04 EF F0 8F EC 13 06 00 01
83 25 C4 FE 13 05 E0 02 EF F0 8F EB 13 06 10 01
83 25 C4 FE 13 05 00 02 EF F0 8F EA 13 06 20 01
83 25 C4 FE 13 05 60 04 EF F0 8F E9 13 06 30 01
83 25 C4 FE 13 05 20 05 EF F0 8F E8 13 06 40 01
83 25 C4 FE 13 05 F0 04 EF F0 8F E7 13 06 50 01
83 25 C4 FE 13 05 D0 04 EF F0 8F E6 13 06 60 01
83 25 C4 FE 13 05 00 02 EF F0 8F E5 13 06 70 01
83 25 C4 FE 13 05 00 02 EF F0 8F E4 13 06 80 01
83 25 C4 FE 13 05 40 05 EF F0 8F E3 13 06 90 01
83 25 C4 FE 13 05 80 04 EF F0 8F E2 13 06 A0 01
83 25 C4 FE 13 05 20 05 EF F0 8F E1 13 06 B0 01
83 25 C4 FE 13 05 50 04 EF F0 8F E0 13 06 C0 01
83 25 C4 FE 13 05 10 04 EF F0 8F DF 13 06 D0 01
83 25 C4 FE 13 05 40 04 EF F0 8F DE 13 06 E0 01
83 25 C4 FE 13 05 00 02 EF F0 8F DD B7 07 C0 00
03 A7 07 00 93 07 40 00 63 1A F7 00 13 06 F0 01
83 25 C4 FE 13 05 00 03 EF F0 8F DB B7 07 C0 00
03 A7 07 00 93 07 50 00 63 1A F7 00 13 06 F0 01
83 25 C4 FE 13 05 10 03 EF F0 8F D9 B7 07 C0 00
03 A7 07 00 93 07 60 00 63 1A F7 00 13 06 F0 01
83 25 C4 FE 13 05 20 03 EF F0 8F D7 B7 07 C0 00
03 A7 07 00 93 07 70 00 63 1A F7 00 13 06 F0 01
83 25 C4 FE 13 05 30 03 EF F0 8F D5 B7 07 C0 00
03 A7 07 00 93 07 80 00 63 1A F7 00 13 06 F0 01
83 25 C4 FE 13 05 40 03 EF F0 8F D3 B7 07 C0 00
03 A7 07 00 93 07 90 00 63 1A F7 00 13 06 F0 01
83 25 C4 FE 13 05 50 03 EF F0 8F D1 B7 07 C0 00
03 A7 07 00 93 07 A0 00 63 1A F7 00 13 06 F0 01
83 25 C4 FE 13 05 60 03 EF F0 8F CF B7 07 C0 00
03 A7 07 00 93 07 B0 00 63 1A F7 00 13 06 F0 01
83 25 C4 FE 13 05 70 03 EF F0 8F CD 13 00 00 00
83 20 C1 01 03 24 81 01 13 01 01 02 67 80 00 00
13 01 01 F9 23 26 11 06 23 24 81 06 13 04 01 07
B7 07 C0 00 93 87 47 00 83 A7 07 00 23 22 F4 FE
B7 07 C0 00 83 A7 07 00 23 20 F4 FE 23 2E 04 FC
93 07 80 04 23 26 F4 FC 93 07 90 04 23 28 F4 FC
23 2A 04 FC 93 07 00 02 23 20 F4 FC 93 07 A0 00
23 22 F4 FC 23 24 04 FC 93 07 10 03 23 2A F4 FA
93 07 A0 00 23 2C F4 FA 23 2E 04 FA 93 07 20 03
23 24 F4 FA 93 07 A0 00 23 26 F4 FA 23 28 04 FA
93 07 30 03 23 2E F4 F8 93 07 A0 00 23 20 F4 FA
23 22 04 FA EF F0 8F E3 23 26 04 FE 6F 00 80 04
23 24 04 FE 6F 00 80 02 B7 17 40 00 93 87 07 80
03 26 C4 FE 83 25 84 FE 13 85 07 00 EF F0 4F C0
83 27 84 FE 93 87 17 00 23 24 F4 FE 03 27 84 FE
93 07 70 00 E3 DA E7 FC 83 27 C4 FE 93 87 17 00
23 26 F4 FE 03 27 84 FD 93 07 E0 01 E3 DA E7 FA
03 27 04 FE 93 07 70 00 63 08 F7 14 03 27 04 FE
93 07 70 00 63 C0 E7 18 03 27 04 FE 93 07 60 00
63 00 F7 0E 03 27 04 FE 93 07 60 00 63 C4 E7 16
03 27 04 FE 93 07 40 00 63 0A F7 00 03 27 04 FE
93 07 50 00 63 00 F7 04 6F 00 C0 14 B7 27 C0 03
93 87 47 02 83 A7 07 00 63 96 07 00 13 05 00 00
EF F0 9F BE B7 27 C0 03 93 87 47 02 03 A7 07 00
93 07 40 00 63 D2 E7 12 13 05 00 00 EF F0 DF BC
6F 00 80 11 B7 27 C0 03 93 87 47 02 03 A7 07 00
93 07 10 00 63 16 F7 00 13 05 20 00 EF F0 DF BA
B7 27 C0 03 93 87 47 02 03 A7 07 00 93 07 40 00
63 D6 E7 00 13 05 20 00 EF F0 1F B9 13 06 00 00
93 05 A0 00 13 05 B0 02 EF F0 8F B0 13 06 10 00
93 05 A0 00 13 05 B0 02 EF F0 8F AF 13 06 20 00
93 05 A0 00 13 05 B0 02 EF F0 8F AE 13 06 30 00
93 05 A0 00 13 05 B0 02 EF F0 8F AD 6F 00 00 00
B7 27 C0 03 93 87 47 02 03 A7 07 00 93 07 20 00
63 16 F7 00 13 05 40 00 EF F0 1F B3 B7 27 C0 03
93 87 47 02 03 A7 07 00 93 07 40 00 63 D6 E7 00
13 05 40 00 EF F0 5F B1 B7 27 C0 03 93 87 47 02
03 A7 07 00 93 07 40 00 63 D6 E7 00 13 05 40 00
EF F0 9F AF 6F 00 00 00 B7 27 C0 03 93 87 47 02
03 A7 07 00 93 07 30 00 63 16 F7 00 13 05 60 00
EF F0 9F AD B7 27 C0 03 93 87 47 02 03 A7 07 00
93 07 40 00 63 D6 E7 00 13 05 60 00 EF F0 DF AB
6F 00 00 00 6F 00 00 00 13 00 00 00 6F F0 5F E6
