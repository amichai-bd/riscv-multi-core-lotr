@00400000
00 00 C0 3F CD CC 0C 40 DC 08 00 00 68 09 00 00
E8 08 00 00 68 09 00 00 58 09 00 00 68 09 00 00
E8 08 00 00 DC 08 00 00 DC 08 00 00 58 09 00 00
E8 08 00 00 B8 08 00 00 B8 08 00 00 B8 08 00 00
F0 08 00 00 00 01 02 02 03 03 03 03 04 04 04 04
04 04 04 04 05 05 05 05 05 05 05 05 05 05 05 05
05 05 05 05 06 06 06 06 06 06 06 06 06 06 06 06
06 06 06 06 06 06 06 06 06 06 06 06 06 06 06 06
06 06 06 06 07 07 07 07 07 07 07 07 07 07 07 07
07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07
07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07
07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07
07 07 07 07 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08
