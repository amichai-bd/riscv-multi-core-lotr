@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 40 38 73 00 10 00
@000000A8
13 01 01 FD 23 26 81 02 13 04 01 03 93 07 05 00
23 2C B4 FC 23 2A C4 FC A3 0F F4 FC 03 27 84 FD
93 07 07 00 93 97 27 00 B3 87 E7 00 93 97 67 00
23 26 F4 FE 83 27 44 FD 93 97 27 00 23 24 F4 FE
03 27 84 FE 83 27 C4 FE 33 07 F7 00 B7 07 40 03
B3 07 F7 00 23 22 F4 FE 03 27 84 FE 83 27 C4 FE
33 07 F7 00 B7 07 40 03 93 87 07 14 B3 07 F7 00
23 20 F4 FE 83 47 F4 FD 37 07 40 00 13 07 87 0A
93 97 27 00 B3 07 F7 00 83 A7 07 00 13 87 07 00
83 27 44 FE 23 A0 E7 00 83 47 F4 FD 37 07 40 00
13 07 C7 22 93 97 27 00 B3 07 F7 00 83 A7 07 00
13 87 07 00 83 27 04 FE 23 A0 E7 00 13 00 00 00
03 24 C1 02 13 01 01 03 67 80 00 00 13 01 01 FD
23 26 11 02 23 24 81 02 13 04 01 03 23 2E A4 FC
23 26 04 FE 23 24 04 FE 23 22 04 FE B7 07 C0 00
93 87 07 22 83 A7 07 00 23 22 F4 FE B7 07 C0 00
93 87 47 23 83 A7 07 00 23 24 F4 FE 6F 00 80 0B
83 27 C4 FE 03 27 C4 FD B3 07 F7 00 03 C7 07 00
93 07 A0 00 63 1A F7 02 23 22 04 FE 83 27 84 FE
93 87 27 00 23 24 F4 FE 03 27 84 FE 93 07 80 07
63 14 F7 00 23 24 04 FE 83 27 C4 FE 93 87 17 00
23 26 F4 FE 6F 00 00 07 83 27 C4 FE 03 27 C4 FD
B3 07 F7 00 83 C7 07 00 03 27 84 FE 83 26 44 FE
13 86 06 00 93 05 07 00 13 85 07 00 EF F0 5F E8
83 27 44 FE 93 87 17 00 23 22 F4 FE 03 27 44 FE
93 07 00 05 63 12 F7 02 23 22 04 FE 83 27 84 FE
93 87 27 00 23 24 F4 FE 03 27 84 FE 93 07 80 07
63 14 F7 00 23 24 04 FE 83 27 C4 FE 93 87 17 00
23 26 F4 FE 83 27 C4 FE 03 27 C4 FD B3 07 F7 00
83 C7 07 00 E3 9E 07 F2 B7 07 C0 00 93 87 07 22
03 27 44 FE 23 A0 E7 00 B7 07 C0 00 93 87 47 23
03 27 84 FE 23 A0 E7 00 13 00 00 00 83 20 C1 02
03 24 81 02 13 01 01 03 67 80 00 00 13 01 01 FD
23 26 81 02 13 04 01 03 23 2E A4 FC 23 2C B4 FC
23 2A C4 FC 03 27 84 FD 93 07 07 00 93 97 27 00
B3 87 E7 00 93 97 67 00 23 26 F4 FE 83 27 44 FD
93 97 27 00 23 24 F4 FE 03 27 84 FE 83 27 C4 FE
33 07 F7 00 B7 07 40 03 B3 07 F7 00 23 22 F4 FE
03 27 84 FE 83 27 C4 FE 33 07 F7 00 B7 07 40 03
93 87 07 14 B3 07 F7 00 23 20 F4 FE B7 07 40 00
13 87 07 3B 83 27 C4 FD 93 97 27 00 B3 07 F7 00
83 A7 07 00 13 87 07 00 83 27 44 FE 23 A0 E7 00
B7 07 40 00 13 87 47 3C 83 27 C4 FD 93 97 27 00
B3 07 F7 00 83 A7 07 00 13 87 07 00 83 27 04 FE
23 A0 E7 00 13 00 00 00 03 24 C1 02 13 01 01 03
67 80 00 00 13 01 01 FE 23 2E 81 00 13 04 01 02
23 26 A4 FE 23 24 B4 FE B7 07 C0 00 93 87 07 22
03 27 84 FE 23 A0 E7 00 B7 07 C0 00 93 87 47 23
03 27 C4 FE 23 A0 E7 00 13 00 00 00 03 24 C1 01
13 01 01 02 67 80 00 00 13 01 01 FE 23 2E 81 00
13 04 01 02 23 26 04 FE B7 07 40 03 23 24 F4 FE
23 26 04 FE 6F 00 40 02 83 27 C4 FE 93 97 27 00
03 27 84 FE B3 07 F7 00 23 A0 07 00 83 27 C4 FE
93 87 17 00 23 26 F4 FE 03 27 C4 FE B7 27 00 00
93 87 F7 57 E3 DA E7 FC 13 00 00 00 13 00 00 00
03 24 C1 01 13 01 01 02 67 80 00 00 13 01 01 FE
23 2E 11 00 23 2C 81 00 13 04 01 02 B7 07 C0 00
83 A7 07 00 23 26 F4 FE 83 27 C4 FE 93 87 C7 FF
13 07 40 00 63 68 F7 10 13 97 27 00 B7 07 40 00
93 87 47 09 B3 07 F7 00 83 A7 07 00 67 80 07 00
B7 07 40 00 13 85 07 00 EF F0 5F D0 13 06 F0 00
93 05 F0 00 13 05 00 00 EF F0 5F E3 13 06 00 01
93 05 F0 00 13 05 10 00 EF F0 5F E2 13 06 10 01
93 05 F0 00 13 05 20 00 EF F0 5F E1 13 06 20 01
93 05 F0 00 13 05 30 00 EF F0 5F E0 13 06 30 01
93 05 F0 00 13 05 40 00 EF F0 5F DF 93 05 00 00
13 05 A0 00 EF F0 1F EB B7 07 40 00 13 85 87 02
EF F0 DF C9 93 05 00 00 13 05 40 01 EF F0 9F E9
B7 07 40 00 13 85 07 05 EF F0 5F C8 93 05 00 00
13 05 E0 01 EF F0 1F E8 B7 07 40 00 13 85 87 08
EF F0 DF C6 13 06 F0 00 93 05 A0 00 13 05 00 00
EF F0 DF D9 13 06 00 01 93 05 A0 00 13 05 10 00
EF F0 DF D8 13 06 10 01 93 05 A0 00 13 05 20 00
EF F0 DF D7 13 06 20 01 93 05 A0 00 13 05 30 00
EF F0 DF D6 13 06 30 01 93 05 A0 00 13 05 40 00
EF F0 DF D5 6F 00 00 00
