@00400800
00 00 C0 3F CD CC 0C 40 EC 08 00 00 78 09 00 00
F8 08 00 00 78 09 00 00 68 09 00 00 78 09 00 00
F8 08 00 00 EC 08 00 00 EC 08 00 00 68 09 00 00
F8 08 00 00 C8 08 00 00 C8 08 00 00 C8 08 00 00
00 09 00 00 D8 0B 00 00 D8 0B 00 00 FC 0B 00 00
D0 0B 00 00 D0 0B 00 00 64 0C 00 00 FC 0B 00 00
D0 0B 00 00 64 0C 00 00 D0 0B 00 00 FC 0B 00 00
CC 0B 00 00 CC 0B 00 00 CC 0B 00 00 64 0C 00 00
00 01 02 02 03 03 03 03 04 04 04 04 04 04 04 04
05 05 05 05 05 05 05 05 05 05 05 05 05 05 05 05
06 06 06 06 06 06 06 06 06 06 06 06 06 06 06 06
06 06 06 06 06 06 06 06 06 06 06 06 06 06 06 06
07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07
07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07
07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07
07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
