@00400000
0C 00 00 00 02 00 00 00 00 00 00 00 06 00 00 00
0A 00 00 00 12 00 00 00 64 00 00 00 04 00 00 00
06 00 00 00 01 00 00 00 00 00 00 00 03 00 00 00
05 00 00 00 09 00 00 00 32 00 00 00 02 00 00 00
1C 02 00 00 68 02 00 00 00 03 00 00 04 03 00 00
08 03 00 00 A0 03 00 00 D4 03 00 00 D8 03 00 00
