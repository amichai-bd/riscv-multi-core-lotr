@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
6F 00 40 06 67 80 00 00
@00000088
13 01 81 FE 23 2A 11 00 23 28 81 00 13 04 81 01
93 07 50 00 23 28 F4 FE 93 07 30 00 23 26 F4 FE
83 25 C4 FE 03 25 04 FF EF 00 40 08 93 07 05 00
23 24 F4 FE B7 17 00 00 93 87 07 F0 03 27 84 FE
23 A0 E7 00 93 07 00 00 13 85 07 00 83 20 41 01
03 24 01 01 13 01 81 01 67 80 00 00 93 00 00 00
13 81 00 00 93 81 00 00 13 82 00 00 93 82 00 00
13 83 00 00 93 83 00 00 13 84 00 00 93 84 00 00
13 85 00 00 93 85 00 00 13 86 00 00 93 86 00 00
13 87 00 00 93 87 00 00 17 11 00 00 13 01 01 DE
13 05 00 00 93 05 00 00 EF F0 9F F5 13 06 05 00
13 05 00 00 93 F6 15 00 63 84 06 00 33 05 C5 00
93 D5 15 00 13 16 16 00 E3 96 05 FE 67 80 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
