@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 C0 43 73 00 10 00
@000000A8
13 01 01 FE 23 2E 81 00 13 04 01 02 23 26 04 FE
6F 00 00 01 83 27 C4 FE 93 87 17 00 23 26 F4 FE
03 27 C4 FE B7 47 01 00 93 87 F7 87 E3 D4 E7 FE
13 00 00 00 13 00 00 00 03 24 C1 01 13 01 01 02
67 80 00 00 13 01 01 FD 23 26 81 02 13 04 01 03
23 2E A4 FC 23 2C B4 FC 23 2A C4 FC 23 28 D4 FC
83 27 84 FD 93 87 17 14 93 97 17 00 03 27 44 FD
B3 07 F7 00 23 22 F4 FE 03 27 C4 FD 93 07 07 00
93 97 27 00 B3 87 E7 00 93 97 47 00 93 87 17 00
23 20 F4 FE 23 26 04 FE 6F 00 40 03 03 27 44 FE
83 27 C4 FE 33 07 F7 40 83 27 04 FD B3 07 F7 00
13 97 27 00 B7 07 40 03 B3 07 F7 00 23 A0 07 00
83 27 C4 FE 93 87 07 05 23 26 F4 FE 03 27 C4 FE
93 07 00 64 E3 D4 E7 FC 23 24 04 FE 6F 00 80 03
03 27 44 FE 83 27 84 FE 33 07 F7 40 83 27 04 FD
B3 07 F7 00 13 97 27 00 B7 07 40 03 B3 07 F7 00
13 07 F0 FF 23 A0 E7 00 83 27 84 FE 93 87 07 05
23 24 F4 FE 03 27 84 FE 83 27 04 FE E3 42 F7 FC
13 00 00 00 13 00 00 00 03 24 C1 02 13 01 01 03
67 80 00 00 13 01 01 FD 23 26 81 02 13 04 01 03
23 2E A4 FC 23 2C B4 FC 83 27 C4 FD 83 A7 07 00
23 26 F4 FE 83 27 84 FD 03 A7 07 00 83 27 C4 FD
23 A0 E7 00 83 27 84 FD 03 27 C4 FE 23 A0 E7 00
13 00 00 00 03 24 C1 02 13 01 01 03 67 80 00 00
13 01 01 FD 23 26 11 02 23 24 81 02 13 04 01 03
23 2E A4 FC 23 2C B4 FC 23 2A C4 FC 23 28 D4 FC
23 26 04 FE 6F 00 C0 0F 23 24 04 FE 6F 00 00 0D
83 27 84 FE 93 97 27 00 03 27 C4 FD B3 07 F7 00
03 A7 07 00 83 27 84 FE 93 87 17 00 93 97 27 00
83 26 C4 FD B3 87 F6 00 83 A7 07 00 63 DA E7 08
83 27 84 FE 93 97 27 00 03 27 C4 FD B3 06 F7 00
83 27 84 FE 93 87 17 00 93 97 27 00 03 27 C4 FD
B3 07 F7 00 93 85 07 00 13 85 06 00 EF F0 9F F2
83 27 84 FE 93 97 27 00 03 27 C4 FD B3 07 F7 00
83 A7 07 00 83 26 04 FD 03 26 44 FD 83 25 84 FE
13 85 07 00 EF F0 1F E1 83 27 84 FE 93 87 17 00
93 97 27 00 03 27 C4 FD B3 07 F7 00 03 A7 07 00
83 27 84 FE 93 87 17 00 83 26 04 FD 03 26 44 FD
93 85 07 00 13 05 07 00 EF F0 DF DD EF F0 5F D9
83 27 84 FE 93 87 17 00 23 24 F4 FE 03 27 84 FD
83 27 C4 FE B3 07 F7 40 93 87 F7 FF 03 27 84 FE
E3 40 F7 F2 83 27 C4 FE 93 87 17 00 23 26 F4 FE
83 27 84 FD 93 87 F7 FF 03 27 C4 FE E3 4E F7 EE
13 00 00 00 13 00 00 00 83 20 C1 02 03 24 81 02
13 01 01 03 67 80 00 00 13 01 01 FD 23 26 11 02
23 24 81 02 13 04 01 03 23 2E A4 FC 23 2C B4 FC
23 2A C4 FC 23 28 D4 FC 93 07 10 00 23 26 F4 FE
6F 00 00 12 83 27 C4 FE 93 97 27 00 03 27 C4 FD
B3 07 F7 00 83 A7 07 00 23 22 F4 FE 83 27 C4 FE
93 87 F7 FF 23 24 F4 FE 6F 00 40 07 83 27 84 FE
93 97 27 00 03 27 C4 FD 33 07 F7 00 83 27 84 FE
93 87 17 00 93 97 27 00 83 26 C4 FD B3 87 F6 00
03 27 07 00 23 A0 E7 00 83 27 84 FE 93 87 17 00
93 97 27 00 03 27 C4 FD B3 07 F7 00 03 A7 07 00
83 27 84 FE 93 87 17 00 83 26 04 FD 03 26 44 FD
93 85 07 00 13 05 07 00 EF F0 DF CC EF F0 5F C8
83 27 84 FE 93 87 F7 FF 23 24 F4 FE 83 27 84 FE
63 C0 07 02 83 27 84 FE 93 97 27 00 03 27 C4 FD
B3 07 F7 00 83 A7 07 00 03 27 44 FE E3 48 F7 F6
83 27 84 FE 93 87 17 00 93 97 27 00 03 27 C4 FD
B3 07 F7 00 03 27 44 FE 23 A0 E7 00 83 27 84 FE
93 87 17 00 93 97 27 00 03 27 C4 FD B3 07 F7 00
03 A7 07 00 83 27 84 FE 93 87 17 00 83 26 04 FD
03 26 44 FD 93 85 07 00 13 05 07 00 EF F0 9F C4
EF F0 1F C0 83 27 C4 FE 93 87 17 00 23 26 F4 FE
03 27 C4 FE 83 27 84 FD E3 4E F7 EC 13 00 00 00
13 00 00 00 83 20 C1 02 03 24 81 02 13 01 01 03
67 80 00 00 13 01 01 F6 23 2E 11 08 23 2C 81 08
13 04 01 0A B7 07 C0 00 83 A7 07 00 23 24 F4 FC
83 27 84 FC 93 87 C7 FF 13 07 70 00 63 64 F7 6A
13 97 27 00 B7 07 40 00 93 87 07 12 B3 07 F7 00
83 A7 07 00 67 80 07 00 EF F0 9F B8 B7 07 40 00
13 87 07 00 93 07 04 F6 93 06 07 00 13 07 80 04
13 06 07 00 93 85 06 00 13 85 07 00 EF 00 C0 66
93 07 20 01 23 24 F4 FA 23 24 04 FE 6F 00 C0 03
83 27 84 FE 93 97 27 00 13 07 04 FF B3 07 F7 00
03 A7 07 F7 B7 17 00 00 93 86 07 E1 13 06 00 00
83 25 84 FE 13 05 07 00 EF F0 DF B6 83 27 84 FE
93 87 17 00 23 24 F4 FE 03 27 84 FE 83 27 84 FA
E3 40 F7 FC EF F0 DF B0 13 07 04 F6 B7 17 00 00
93 86 07 E1 13 06 00 00 83 25 84 FA 13 05 07 00
EF F0 1F C7 EF F0 DF AE 6F F0 1F F6 EF F0 5F AE
B7 07 40 00 13 87 87 04 93 07 04 F6 93 06 07 00
13 07 80 04 13 06 07 00 93 85 06 00 13 85 07 00
EF 00 80 5C 93 07 20 01 23 26 F4 FA 23 22 04 FE
6F 00 00 04 83 27 44 FE 93 97 27 00 13 07 04 FF
B3 07 F7 00 03 A7 07 F7 B7 17 00 00 93 86 07 E1
B7 17 00 00 13 86 87 2E 83 25 44 FE 13 05 07 00
EF F0 5F AC 83 27 44 FE 93 87 17 00 23 22 F4 FE
03 27 44 FE 83 27 C4 FA E3 4E F7 FA EF F0 5F A6
13 07 04 F6 B7 17 00 00 93 86 07 E1 B7 17 00 00
13 86 87 2E 83 25 C4 FA 13 05 07 00 EF F0 5F BC
EF F0 1F A4 6F F0 9F F5 23 26 04 FE 6F 00 C0 0B
83 27 C4 FE 13 97 27 00 B7 07 40 03 B3 07 F7 00
13 07 F0 FF 23 A0 E7 00 03 27 C4 FE B7 17 00 00
93 87 07 96 B3 07 F7 00 13 97 27 00 B7 07 40 03
93 87 07 EC B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
03 27 C4 FE B7 17 00 00 93 87 07 2C B3 07 F7 00
13 97 27 00 B7 07 40 03 93 87 07 EC B3 07 F7 00
13 07 F0 FF 23 A0 E7 00 03 27 C4 FE B7 27 00 00
93 87 07 C2 B3 07 F7 00 13 97 27 00 B7 07 40 03
93 87 07 EC B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
83 27 C4 FE 13 97 27 00 B7 97 40 03 93 87 07 4C
B3 07 F7 00 13 07 F0 FF 23 A0 E7 00 83 27 C4 FE
93 87 17 00 23 26 F4 FE 03 27 C4 FE 93 07 F0 04
E3 D0 E7 F4 23 26 04 FE 6F 00 00 09 03 27 C4 FE
93 07 07 00 93 97 27 00 B3 87 E7 00 93 97 67 00
13 87 07 00 B7 07 40 03 B3 07 F7 00 13 07 F0 FF
23 A0 E7 00 03 27 C4 FE 93 07 07 00 93 97 27 00
B3 87 E7 00 93 97 67 00 13 87 07 00 B7 07 40 03
93 87 C7 09 B3 07 F7 00 13 07 F0 FF 23 A0 E7 00
03 27 C4 FE 93 07 07 00 93 97 27 00 B3 87 E7 00
93 97 67 00 13 87 07 00 B7 07 40 03 93 87 C7 13
B3 07 F7 00 13 07 F0 FF 23 A0 E7 00 83 27 C4 FE
93 87 17 00 23 26 F4 FE 03 27 C4 FE 93 07 70 07
E3 D6 E7 F6 EF F0 DF 8C B7 07 40 00 13 87 07 09
93 07 04 F6 93 06 07 00 13 07 80 04 13 06 07 00
93 85 06 00 13 85 07 00 EF 00 00 3B 93 07 20 01
23 28 F4 FA 23 20 04 FE 6F 00 C0 03 83 27 04 FE
93 97 27 00 13 07 04 FF B3 07 F7 00 03 A7 07 F7
B7 17 00 00 93 86 07 E1 13 06 80 02 83 25 04 FE
13 05 07 00 EF F0 1F 8B 83 27 04 FE 93 87 17 00
23 20 F4 FE 03 27 04 FE 83 27 04 FB E3 40 F7 FC
EF F0 1F 85 13 07 04 F6 B7 17 00 00 93 86 07 E1
13 06 80 02 83 25 04 FB 13 05 07 00 EF F0 5F 9B
EF F0 1F 83 6F F0 1F F6 EF F0 9F 82 B7 07 40 00
13 87 87 0D 93 07 04 F6 93 06 07 00 13 07 80 04
13 06 07 00 93 85 06 00 13 85 07 00 EF 00 C0 30
93 07 20 01 23 2A F4 FA 23 2E 04 FC 6F 00 00 04
83 27 C4 FD 93 97 27 00 13 07 04 FF B3 07 F7 00
03 A7 07 F7 B7 17 00 00 93 86 07 E1 B7 17 00 00
13 86 07 2C 83 25 C4 FD 13 05 07 00 EF F0 9F 80
83 27 C4 FD 93 87 17 00 23 2E F4 FC 03 27 C4 FD
83 27 44 FB E3 4E F7 FA EF F0 8F FA 13 07 04 F6
B7 17 00 00 93 86 07 E1 B7 17 00 00 13 86 07 2C
83 25 44 FB 13 05 07 00 EF F0 9F 90 EF F0 4F F8
6F F0 9F F5 EF F0 CF F7 B7 07 40 00 13 87 07 00
93 07 04 F6 93 06 07 00 13 07 80 04 13 06 07 00
93 85 06 00 13 85 07 00 EF 00 00 26 93 07 20 01
23 2C F4 FA 23 2C 04 FC 6F 00 80 03 83 27 84 FD
93 97 27 00 13 07 04 FF B3 07 F7 00 83 A7 07 F7
93 06 00 4B 13 06 00 00 83 25 84 FD 13 85 07 00
EF F0 4F F6 83 27 84 FD 93 87 17 00 23 2C F4 FC
03 27 84 FD 83 27 84 FB E3 42 F7 FC EF F0 4F F0
93 07 04 F6 93 06 00 4B 13 06 00 00 83 25 84 FB
13 85 07 00 EF F0 5F 9B EF F0 8F EE 6F F0 9F F6
EF F0 0F EE B7 07 40 00 13 87 87 04 93 07 04 F6
93 06 07 00 13 07 80 04 13 06 07 00 93 85 06 00
13 85 07 00 EF 00 40 1C 93 07 20 01 23 2E F4 FA
23 2A 04 FC 6F 00 C0 03 83 27 44 FD 93 97 27 00
13 07 04 FF B3 07 F7 00 03 A7 07 F7 93 06 00 4B
B7 17 00 00 13 86 87 2E 83 25 44 FD 13 05 07 00
EF F0 4F EC 83 27 44 FD 93 87 17 00 23 2A F4 FC
03 27 44 FD 83 27 C4 FB E3 40 F7 FC EF F0 4F E6
13 07 04 F6 93 06 00 4B B7 17 00 00 13 86 87 2E
83 25 C4 FB 13 05 07 00 EF F0 1F 91 EF F0 4F E4
6F F0 1F F6 EF F0 CF E3 B7 07 40 00 13 87 07 09
93 07 04 F6 93 06 07 00 13 07 80 04 13 06 07 00
93 85 06 00 13 85 07 00 EF 00 00 12 93 07 20 01
23 20 F4 FC 23 28 04 FC 6F 00 80 03 83 27 04 FD
93 97 27 00 13 07 04 FF B3 07 F7 00 83 A7 07 F7
93 06 00 4B 13 06 80 02 83 25 04 FD 13 85 07 00
EF F0 4F E2 83 27 04 FD 93 87 17 00 23 28 F4 FC
03 27 04 FD 83 27 04 FC E3 42 F7 FC EF F0 4F DC
93 07 04 F6 93 06 00 4B 13 06 80 02 83 25 04 FC
13 85 07 00 EF F0 5F 87 EF F0 8F DA 6F F0 9F F6
EF F0 0F DA B7 07 40 00 13 87 87 0D 93 07 04 F6
93 06 07 00 13 07 80 04 13 06 07 00 93 85 06 00
13 85 07 00 EF 00 40 08 93 07 20 01 23 22 F4 FC
23 26 04 FC 6F 00 C0 03 83 27 C4 FC 93 97 27 00
13 07 04 FF B3 07 F7 00 03 A7 07 F7 93 06 00 4B
B7 17 00 00 13 86 07 2C 83 25 C4 FC 13 05 07 00
EF F0 4F D8 83 27 C4 FC 93 87 17 00 23 26 F4 FC
03 27 C4 FC 83 27 44 FC E3 40 F7 FC EF F0 4F D2
13 07 04 F6 93 06 00 4B B7 17 00 00 13 86 07 2C
83 25 44 FC 13 05 07 00 EF F0 0F FD EF F0 4F D0
6F F0 1F F6 6F 00 00 00 B3 C7 A5 00 93 F7 37 00
B3 08 C5 00 63 96 07 06 93 07 30 00 63 F2 C7 06
93 77 35 00 13 07 05 00 63 9A 07 0C 13 F6 C8 FF
B3 06 E6 40 93 07 00 02 93 02 00 02 63 C2 D7 06
93 86 05 00 93 07 07 00 63 78 C7 02 03 A8 06 00
93 87 47 00 93 86 46 00 23 AE 07 FF E3 E8 C7 FE
93 07 F6 FF B3 87 E7 40 93 F7 C7 FF 93 87 47 00
33 07 F7 00 B3 85 F5 00 63 68 17 01 67 80 00 00
13 07 05 00 E3 7C 15 FF 83 C7 05 00 13 07 17 00
93 85 15 00 A3 0F F7 FE E3 68 17 FF 67 80 00 00
83 A6 45 00 83 A7 C5 01 83 AF 05 00 03 AF 85 00
83 AE C5 00 03 AE 05 01 03 A3 45 01 03 A8 85 01
23 22 D7 00 83 A6 05 02 23 20 F7 01 23 24 E7 01
23 26 D7 01 23 28 C7 01 23 2A 67 00 23 2C 07 01
23 2E F7 00 13 07 47 02 B3 07 E6 40 23 2E D7 FE
93 85 45 02 E3 C6 F2 FA 6F F0 9F F4 83 C6 05 00
13 07 17 00 93 77 37 00 A3 0F D7 FE 93 85 15 00
E3 8E 07 F0 83 C6 05 00 13 07 17 00 93 77 37 00
A3 0F D7 FE 93 85 15 00 E3 9A 07 FC 6F F0 1F F0
