@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 C0 21
@00000018
13 01 01 FE 23 2E 11 00 23 2C 81 00 13 04 01 02
93 07 40 01 23 26 F4 FE 93 07 50 00 23 24 F4 FE
83 25 84 FE 03 25 C4 FE EF 00 C0 23 93 07 05 00
23 22 F4 FE 83 27 44 FE 13 85 07 00 83 20 C1 01
03 24 81 01 13 01 01 02 67 80 00 00 13 01 01 FE
23 2E 11 00 23 2C 81 00 13 04 01 02 93 07 80 00
23 26 F4 FE 93 07 90 01 23 24 F4 FE 83 25 84 FE
03 25 C4 FE EF 00 00 1F 93 07 05 00 23 22 F4 FE
83 27 44 FE 13 85 07 00 83 20 C1 01 03 24 81 01
13 01 01 02 67 80 00 00 13 01 01 FE 23 2E 11 00
23 2C 81 00 13 04 01 02 93 07 A0 00 23 26 F4 FE
93 07 E0 01 23 24 F4 FE 83 25 84 FE 03 25 C4 FE
EF 00 40 1A 93 07 05 00 23 22 F4 FE 83 27 44 FE
13 85 07 00 83 20 C1 01 03 24 81 01 13 01 01 02
67 80 00 00 13 01 01 FE 23 2E 11 00 23 2C 81 00
13 04 01 02 93 07 40 06 23 26 F4 FE 93 07 40 00
23 24 F4 FE 83 25 84 FE 03 25 C4 FE EF 00 80 15
93 07 05 00 23 22 F4 FE 83 27 44 FE 13 85 07 00
83 20 C1 01 03 24 81 01 13 01 01 02 67 80 00 00
13 01 01 FE 23 2E 11 00 23 2C 81 00 23 2A 91 00
13 04 01 02 B7 07 C0 00 93 87 47 00 83 A7 07 00
23 26 F4 FE 03 27 C4 FE 93 07 30 00 63 04 F7 08
03 27 C4 FE 93 07 30 00 63 CA E7 08 03 27 C4 FE
93 07 20 00 63 0C F7 04 03 27 C4 FE 93 07 20 00
63 CE E7 06 83 27 C4 FE 63 8A 07 00 03 27 C4 FE
93 07 10 00 63 00 F7 02 6F 00 40 06 B7 17 40 00
93 84 07 F0 EF F0 DF E5 93 07 05 00 23 A0 F4 00
6F 00 C0 04 B7 17 40 00 93 84 47 F0 EF F0 1F E9
93 07 05 00 23 A0 F4 00 6F 00 40 03 B7 17 40 00
93 84 87 F0 EF F0 5F EC 93 07 05 00 23 A0 F4 00
6F 00 C0 01 B7 17 40 00 93 84 C7 F0 EF F0 9F EF
93 07 05 00 23 A0 F4 00 13 00 00 00 13 00 00 00
13 85 07 00 83 20 C1 01 03 24 81 01 83 24 41 01
13 01 01 02 67 80 00 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF F0 1F ED 13 06 05 00 13 05 00 00 93 F6 15 00
63 84 06 00 33 05 C5 00 93 D5 15 00 13 16 16 00
E3 96 05 FE 67 80 00 00
