@00400800
48 00 00 00 45 00 00 00 4C 00 00 00 4C 00 00 00
4F 00 00 00 20 00 00 00 50 00 00 00 52 00 00 00
49 00 00 00 4E 00 00 00 54 00 00 00 2C 00 00 00
0A 00 00 00 00 00 00 00 30 00 00 00 0A 00 00 00
00 00 00 00 31 00 00 00 0A 00 00 00 00 00 00 00
32 00 00 00 0A 00 00 00 00 00 00 00 33 00 00 00
0A 00 00 00 00 00 00 00
