@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 80 00 73 00 10 00
@000000A8
13 01 01 FB 23 26 81 04 13 04 01 05 B7 07 C0 00
83 A7 07 00 23 28 F4 FC 93 07 10 00 23 26 F4 FE
23 24 04 FE 93 07 F0 3F 23 22 F4 FE 23 26 04 FC
23 20 04 FE 93 07 10 00 23 2E F4 FC 93 07 00 20
23 2C F4 FC 23 2A 04 FC 93 07 E0 07 23 2A F4 FA
93 07 D0 07 23 2C F4 FA 93 07 B0 07 23 2E F4 FA
93 07 70 07 23 20 F4 FC 93 07 F0 06 23 22 F4 FC
93 07 F0 05 23 24 F4 FC 03 27 04 FD 93 07 40 00
63 0A F7 00 03 27 04 FD 93 07 80 00 63 04 F7 34
6F 00 40 3D B7 27 00 03 93 87 47 02 83 A7 07 00
63 9C 07 06 93 07 10 00 23 26 F4 FE 93 07 F0 3F
23 22 F4 FE 23 26 04 FC 93 07 10 00 23 2E F4 FC
93 07 00 20 23 2C F4 FC 6F 00 00 01 83 27 84 FE
93 87 17 00 23 24 F4 FE 03 27 84 FE 93 07 10 68
E3 D6 E7 FE B7 27 00 03 93 87 87 01 03 27 04 FE
23 A0 E7 00 03 27 04 FE 93 07 F0 3F 63 16 F7 00
23 20 04 FE 6F 00 C0 00 93 07 F0 3F 23 20 F4 FE
23 24 04 FE 6F F0 1F F8 B7 27 00 03 93 87 47 02
03 A7 07 00 93 07 10 00 63 1C F7 06 93 07 F0 3F
23 22 F4 FE 23 26 04 FC 23 20 04 FE 93 07 10 00
23 2E F4 FC 93 07 00 20 23 2C F4 FC 6F 00 00 01
83 27 84 FE 93 87 17 00 23 24 F4 FE 03 27 84 FE
93 07 10 68 E3 D6 E7 FE B7 27 00 03 93 87 87 01
03 27 C4 FE 23 A0 E7 00 83 27 C4 FE 93 87 17 00
23 26 F4 FE 03 27 C4 FE 93 07 F0 3F 63 16 F7 00
93 07 10 00 23 26 F4 FE 23 24 04 FE 6F F0 9F EF
B7 27 00 03 93 87 47 02 03 A7 07 00 93 07 20 00
63 1C F7 06 93 07 10 00 23 26 F4 FE 93 07 F0 3F
23 22 F4 FE 23 26 04 FC 23 20 04 FE 93 07 00 20
23 2C F4 FC 6F 00 00 01 83 27 84 FE 93 87 17 00
23 24 F4 FE 03 27 84 FE 93 07 10 68 E3 D6 E7 FE
B7 27 00 03 93 87 87 01 03 27 C4 FD 23 A0 E7 00
83 27 C4 FD 93 97 17 00 23 2E F4 FC 03 27 C4 FD
93 07 00 20 63 D6 E7 00 93 07 10 00 23 2E F4 FC
23 24 04 FE 6F F0 1F E7 B7 27 00 03 93 87 47 02
03 A7 07 00 93 07 30 00 63 1A F7 06 93 07 10 00
23 26 F4 FE 23 26 04 FC 23 20 04 FE 93 07 10 00
23 2E F4 FC 93 07 00 20 23 2C F4 FC 6F 00 00 01
83 27 84 FE 93 87 17 00 23 24 F4 FE 03 27 84 FE
93 07 10 68 E3 D6 E7 FE B7 27 00 03 93 87 87 01
03 27 44 FE 23 A0 E7 00 83 27 44 FE 93 87 F7 FF
23 22 F4 FE 83 27 44 FE 63 96 07 00 93 07 F0 3F
23 22 F4 FE 23 24 04 FE 6F F0 DF DE B7 27 00 03
93 87 47 02 03 A7 07 00 93 07 40 00 63 1E F7 06
93 07 10 00 23 26 F4 FE 93 07 F0 3F 23 22 F4 FE
23 26 04 FC 23 20 04 FE 93 07 10 00 23 2E F4 FC
6F 00 00 01 83 27 84 FE 93 87 17 00 23 24 F4 FE
03 27 84 FE 93 07 10 68 E3 D6 E7 FE B7 27 00 03
93 87 87 01 03 27 84 FD 23 A0 E7 00 83 27 84 FD
13 D7 F7 01 B3 07 F7 00 93 D7 17 40 23 2C F4 FC
83 27 84 FD 63 96 07 00 93 07 00 20 23 2C F4 FC
23 24 04 FE 6F F0 1F D6 B7 27 00 03 93 87 47 02
03 A7 07 00 93 07 50 00 E3 16 F7 D4 93 07 10 00
23 26 F4 FE 93 07 F0 3F 23 22 F4 FE 23 20 04 FE
93 07 10 00 23 2E F4 FC 93 07 00 20 23 2C F4 FC
6F 00 00 01 83 27 84 FE 93 87 17 00 23 24 F4 FE
03 27 84 FE 93 07 30 1F E3 D6 E7 FE 83 27 44 FD
13 87 17 00 23 2A E4 FC 37 27 00 03 93 97 27 00
93 06 04 FF B3 87 F6 00 83 A7 47 FC 23 20 F7 00
03 27 44 FD 93 07 50 00 63 D4 E7 00 23 2A 04 FC
23 24 04 FE 6F F0 1F CD 83 27 84 FE 93 87 17 00
23 24 F4 FE 03 27 84 FE 93 07 90 0F E3 D6 E7 FE
B7 27 00 03 13 87 47 00 83 27 44 FD 93 97 27 00
93 06 04 FF B3 87 F6 00 83 A7 47 FC 23 20 F7 00
B7 27 00 03 13 87 87 00 83 27 44 FD 93 97 27 00
93 06 04 FF B3 87 F6 00 83 A7 47 FC 23 20 F7 00
B7 27 00 03 13 87 C7 00 83 27 44 FD 93 97 27 00
93 06 04 FF B3 87 F6 00 83 A7 47 FC 23 20 F7 00
83 27 44 FD 93 87 17 00 23 2A F4 FC 03 27 44 FD
93 07 50 00 63 D4 E7 00 23 2A 04 FC 23 24 04 FE
6F F0 5F F7 6F 00 00 00
