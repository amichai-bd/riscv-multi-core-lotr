@00400000
03 00 00 00 02 00 00 00 01 00 00 00 04 00 00 00
