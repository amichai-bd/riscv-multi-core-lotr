@00400000
