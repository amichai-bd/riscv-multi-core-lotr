/*
 User handshake FSM 
 Wishbone master unit to 
 handle user handshake 
 between uart host(PC) and lotr
 */

`timescale 1ns/1ns

module handshake
  #()
   (
    input logic clk,
    input logic rstn,
    wishbone.master wb_master
    );

endmodule // handshake

   
