@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 80 00 73 00 10 00
@000000A8
13 01 01 FD 23 26 81 02 13 04 01 03 B7 07 C0 00
93 87 47 00 83 A7 07 00 23 26 F4 FE 93 07 90 00
23 24 F4 FE 93 07 80 00 23 22 F4 FE 93 07 70 00
23 20 F4 FE 93 07 30 01 23 2E F4 FC 03 27 C4 FE
93 07 30 00 63 08 F7 14 03 27 C4 FE 93 07 30 00
63 C0 E7 16 03 27 C4 FE 93 07 20 00 63 0E F7 10
03 27 C4 FE 93 07 20 00 63 C4 E7 14 83 27 C4 FE
63 8A 07 00 03 27 C4 FE 93 07 10 00 63 00 F7 0E
6F 00 00 13 B7 07 C0 00 93 87 87 00 03 A7 07 00
93 07 10 00 63 1E F7 04 93 07 80 0C 23 2C F4 FC
B7 07 C0 02 93 87 07 20 03 27 84 FD 23 A0 E7 00
B7 07 C0 02 93 87 47 20 13 07 10 00 23 A0 E7 00
13 00 00 00 B7 07 C0 01 93 87 47 20 83 A7 07 00
E3 8A 07 FE B7 07 C0 01 13 87 07 20 B7 17 40 00
93 87 07 F0 03 27 07 00 23 A0 E7 00 6F 00 00 07
B7 07 C0 00 93 87 87 00 03 A7 07 00 93 07 20 00
63 1E F7 04 93 07 80 25 23 2C F4 FC B7 07 C0 01
93 87 07 20 03 27 84 FD 23 A0 E7 00 B7 07 C0 01
93 87 47 20 13 07 10 00 23 A0 E7 00 13 00 00 00
B7 07 C0 02 93 87 47 20 83 A7 07 00 E3 8A 07 FE
B7 07 C0 02 13 87 07 20 B7 17 40 00 93 87 07 F0
03 27 07 00 23 A0 E7 00 6F 00 00 00 B7 07 C0 00
93 87 47 15 23 A0 07 00 13 00 00 00 13 00 00 00
23 2C F4 FC 6F 00 C0 03 B7 07 C0 00 93 87 87 15
23 A0 07 00 13 00 00 00 13 00 00 00 23 2C F4 FC
6F 00 00 02 B7 07 C0 00 93 87 C7 15 23 A0 07 00
13 00 00 00 13 00 00 00 23 2C F4 FC 13 00 00 00
93 07 00 00 13 85 07 00 03 24 C1 02 13 01 01 03
67 80 00 00
