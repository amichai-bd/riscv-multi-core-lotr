@00400000
42 55 42 42 4C 45 20 53 4F 52 54 20 52 41 4E 44
4F 4D 0A 00 42 55 42 42 4C 45 20 53 4F 52 54 20
33 20 55 4E 49 51 55 45 0A 00 00 00 42 55 42 42
4C 45 20 53 4F 52 54 20 52 45 56 45 52 53 45 0A
00 00 00 00 42 55 42 42 4C 45 20 53 4F 52 54 20
41 4C 4D 4F 53 54 20 53 4F 52 54 45 44 0A 00 00
49 4E 53 45 52 54 49 4F 4E 20 53 4F 52 54 20 52
41 4E 44 4F 4D 0A 00 00 49 4E 53 45 52 54 49 4F
4E 20 53 4F 52 54 20 33 20 55 4E 49 51 55 45 0A
00 00 00 00 49 4E 53 45 52 54 49 4F 4E 20 53 4F
52 54 20 52 45 56 45 52 53 45 0A 00 49 4E 53 45
52 54 49 4F 4E 20 53 4F 52 54 20 41 4C 4D 4F 53
54 20 53 4F 52 54 45 44 2E 0A 00 00 0B 00 00 00
05 00 00 00 09 00 00 00 0D 00 00 00 12 00 00 00
07 00 00 00 01 00 00 00 02 00 00 00 0C 00 00 00
0A 00 00 00 04 00 00 00 03 00 00 00 0E 00 00 00
06 00 00 00 0F 00 00 00 11 00 00 00 08 00 00 00
10 00 00 00 06 00 00 00 12 00 00 00 0C 00 00 00
0C 00 00 00 06 00 00 00 12 00 00 00 12 00 00 00
06 00 00 00 06 00 00 00 0C 00 00 00 0C 00 00 00
12 00 00 00 06 00 00 00 12 00 00 00 06 00 00 00
0C 00 00 00 12 00 00 00 0C 00 00 00 12 00 00 00
11 00 00 00 10 00 00 00 0F 00 00 00 0E 00 00 00
0D 00 00 00 0C 00 00 00 0B 00 00 00 0A 00 00 00
09 00 00 00 08 00 00 00 07 00 00 00 06 00 00 00
05 00 00 00 04 00 00 00 03 00 00 00 02 00 00 00
01 00 00 00 02 00 00 00 03 00 00 00 04 00 00 00
05 00 00 00 06 00 00 00 07 00 00 00 08 00 00 00
09 00 00 00 0A 00 00 00 0B 00 00 00 0C 00 00 00
0D 00 00 00 0E 00 00 00 0F 00 00 00 10 00 00 00
11 00 00 00 12 00 00 00 01 00 00 00 9C 0A 00 00
58 0B 00 00 1C 0C 00 00 44 0E 00 00 0C 0F 00 00
C0 0F 00 00 7C 10 00 00 30 11 00 00
@0040020C
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 3C 62 52 00 18 1C 1A 00 3C 42 40 00 3C 42 40
00 30 28 24 00 7E 02 3E 00 3C 42 02 00 7E 40 30
00 3C 42 42 00 3C 42 42 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 18 3C 66 00 1E 22 3E 00 3C 3E 02
00 1E 3E 22 00 7E 06 06 00 7E 06 06 00 3C 3E 02
00 66 66 66 00 7E 18 18 00 60 60 60 00 46 66 3E
00 06 06 06 00 42 66 5A 00 62 66 6E 00 3C 66 66
00 3E 66 66 00 3C 42 42 00 3E 66 66 00 7C 06 1E
00 7E 18 18 00 66 66 66 00 66 66 66 00 42 42 42
00 66 66 3C 00 66 66 3C 00 7E 20 10 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 18 18 1E 06 00 00 00 00 00 18 18 00
00 00 00 00 4A 46 3C 00 18 18 7E 00 3C 02 7E 00
38 42 3C 00 7E 20 20 00 40 42 3C 00 3E 42 3C 00
08 08 08 00 3C 42 3C 00 7C 40 3E 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 66 7E 66 00 3E 22 1E 00
02 3E 3C 00 22 3E 1E 00 7E 06 7E 00 7E 06 06 00
3A 22 3C 00 7E 66 66 00 18 18 7E 00 66 66 7C 00
3E 66 46 00 06 06 7E 00 5A 42 42 00 76 66 46 00
66 66 3C 00 3E 06 06 00 52 62 7C 00 3E 66 66 00
78 60 3E 00 18 18 18 00 66 7E 3C 00 66 3C 18 00
5A 7E 42 00 3C 66 66 00 18 18 18 00 08 04 7E 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 30 10 38 7C 30 10 38 38
30 10 38 38 30 10 38 7C 30 10 38 38 00 00 00 00
BA 48 84 82 78 AC 48 44 78 28 28 10 BA 38 10 28
7C 38 48 48 00 00 00 00
