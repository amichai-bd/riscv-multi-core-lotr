@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 80 00 73 00 10 00
@000000A8
13 01 01 FE 23 2E 81 00 13 04 01 02 B7 07 C0 00
93 87 47 00 83 A7 07 00 23 24 F4 FE B7 07 C0 00
83 A7 07 00 23 22 F4 FE 23 26 04 FE 83 27 44 FE
93 87 C7 FF 13 07 70 00 63 6E F7 06 13 97 27 00
B7 17 40 00 93 87 07 80 B3 07 F7 00 83 A7 07 00
67 80 07 00 B7 17 40 02 93 87 07 90 13 07 10 05
23 A0 E7 00 13 00 00 00 83 27 C4 FE 13 87 17 00
23 26 E4 FE 13 07 90 00 E3 58 F7 FE B7 17 40 02
13 87 07 90 B7 17 40 00 93 87 07 F0 03 27 07 00
23 A0 E7 00 6F 00 00 02 6F 00 00 00 6F 00 00 00
6F 00 00 00 6F 00 00 00 6F 00 00 00 6F 00 00 00
6F 00 00 00 93 07 00 00 13 85 07 00 03 24 C1 01
13 01 01 02 67 80 00 00
