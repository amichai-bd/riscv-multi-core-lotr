@00400000
FC 00 00 00 40 01 00 00 44 01 00 00 48 01 00 00
4C 01 00 00 50 01 00 00 54 01 00 00 58 01 00 00
