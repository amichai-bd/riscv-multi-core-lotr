@00400000
00 00 00 00 01 00 00 00 02 00 00 00 03 00 00 00
04 00 00 00 05 00 00 00 06 00 00 00 07 00 00 00
08 00 00 00 09 00 00 00 0A 00 00 00 0B 00 00 00
0C 00 00 00 0D 00 00 00 0E 00 00 00 0F 00 00 00
10 00 00 00 11 00 00 00 12 00 00 00 13 00 00 00
14 00 00 00 15 00 00 00 16 00 00 00 17 00 00 00
18 00 00 00 19 00 00 00 1A 00 00 00 1B 00 00 00
1C 00 00 00 1D 00 00 00 1E 00 00 00 1F 00 00 00
20 00 00 00 21 00 00 00 22 00 00 00 23 00 00 00
24 00 00 00 25 00 00 00 26 00 00 00 27 00 00 00
28 00 00 00 29 00 00 00 2A 00 00 00 2B 00 00 00
2C 00 00 00 2D 00 00 00 2E 00 00 00 2F 00 00 00
30 00 00 00 31 00 00 00 32 00 00 00 33 00 00 00
34 00 00 00 35 00 00 00 36 00 00 00 37 00 00 00
38 00 00 00 39 00 00 00 3A 00 00 00 3B 00 00 00
3C 00 00 00 3D 00 00 00 3E 00 00 00 3F 00 00 00
40 00 00 00 41 00 00 00 42 00 00 00 43 00 00 00
44 00 00 00 45 00 00 00 46 00 00 00 47 00 00 00
48 00 00 00 49 00 00 00 4A 00 00 00 4B 00 00 00
4C 00 00 00 4D 00 00 00 4E 00 00 00 4F 00 00 00
50 00 00 00 51 00 00 00 52 00 00 00 53 00 00 00
54 00 00 00 55 00 00 00 56 00 00 00 57 00 00 00
58 00 00 00 59 00 00 00 5A 00 00 00 5B 00 00 00
5C 00 00 00 5D 00 00 00 5E 00 00 00 5F 00 00 00
60 00 00 00 61 00 00 00 62 00 00 00 63 00 00 00
64 00 00 00 65 00 00 00 66 00 00 00 67 00 00 00
68 00 00 00 69 00 00 00 6A 00 00 00 6B 00 00 00
6C 00 00 00 6D 00 00 00 6E 00 00 00 6F 00 00 00
70 00 00 00 71 00 00 00 72 00 00 00 73 00 00 00
74 00 00 00 75 00 00 00 76 00 00 00 77 00 00 00
78 00 00 00 79 00 00 00 7A 00 00 00 7B 00 00 00
7C 00 00 00 7D 00 00 00 7E 00 00 00 7F 00 00 00
80 00 00 00 81 00 00 00 82 00 00 00 83 00 00 00
84 00 00 00 85 00 00 00 86 00 00 00 87 00 00 00
88 00 00 00 89 00 00 00 8A 00 00 00 8B 00 00 00
8C 00 00 00 8D 00 00 00 8E 00 00 00 8F 00 00 00
8F 00 00 00 8E 00 00 00 8D 00 00 00 8C 00 00 00
8B 00 00 00 8A 00 00 00 89 00 00 00 88 00 00 00
87 00 00 00 86 00 00 00 85 00 00 00 84 00 00 00
83 00 00 00 82 00 00 00 81 00 00 00 80 00 00 00
7F 00 00 00 7E 00 00 00 7D 00 00 00 7C 00 00 00
7B 00 00 00 7A 00 00 00 79 00 00 00 78 00 00 00
77 00 00 00 76 00 00 00 75 00 00 00 74 00 00 00
73 00 00 00 72 00 00 00 71 00 00 00 70 00 00 00
6F 00 00 00 6E 00 00 00 6D 00 00 00 6C 00 00 00
6B 00 00 00 6A 00 00 00 69 00 00 00 68 00 00 00
67 00 00 00 66 00 00 00 65 00 00 00 64 00 00 00
63 00 00 00 62 00 00 00 61 00 00 00 60 00 00 00
5F 00 00 00 5E 00 00 00 5D 00 00 00 5C 00 00 00
5B 00 00 00 5A 00 00 00 59 00 00 00 58 00 00 00
57 00 00 00 56 00 00 00 55 00 00 00 54 00 00 00
53 00 00 00 52 00 00 00 51 00 00 00 50 00 00 00
4F 00 00 00 4E 00 00 00 4D 00 00 00 4C 00 00 00
4B 00 00 00 4A 00 00 00 49 00 00 00 48 00 00 00
47 00 00 00 46 00 00 00 45 00 00 00 44 00 00 00
43 00 00 00 42 00 00 00 41 00 00 00 40 00 00 00
3F 00 00 00 3E 00 00 00 3D 00 00 00 3C 00 00 00
3B 00 00 00 3A 00 00 00 39 00 00 00 38 00 00 00
37 00 00 00 36 00 00 00 35 00 00 00 34 00 00 00
33 00 00 00 32 00 00 00 31 00 00 00 30 00 00 00
2F 00 00 00 2E 00 00 00 2D 00 00 00 2C 00 00 00
2B 00 00 00 2A 00 00 00 29 00 00 00 28 00 00 00
27 00 00 00 26 00 00 00 25 00 00 00 24 00 00 00
23 00 00 00 22 00 00 00 21 00 00 00 20 00 00 00
1F 00 00 00 1E 00 00 00 1D 00 00 00 1C 00 00 00
1B 00 00 00 1A 00 00 00 19 00 00 00 18 00 00 00
17 00 00 00 16 00 00 00 15 00 00 00 14 00 00 00
13 00 00 00 12 00 00 00 11 00 00 00 10 00 00 00
0F 00 00 00 0E 00 00 00 0D 00 00 00 0C 00 00 00
0B 00 00 00 0A 00 00 00 09 00 00 00 08 00 00 00
07 00 00 00 06 00 00 00 05 00 00 00 04 00 00 00
03 00 00 00 02 00 00 00 01 00 00 00 00 00 00 00
