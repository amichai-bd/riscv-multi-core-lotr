`timescale 1ns/1ns

`include "lotr_defines.sv"
module uart_io_tb ();
import lotr_pkg::*;

endmodule