@00400000
02 00 00 00 03 00 00 00 04 00 00 00 0A 00 00 00
28 00 00 00
