@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
6F 00 00 69 67 80 00 00
@00000088
13 01 01 FE 23 2E 81 00 13 04 01 02 23 26 A4 FE
B7 17 40 00 93 87 07 80 03 27 C4 FE 13 07 17 00
23 A0 E7 00 13 00 00 00 03 24 C1 01 13 01 01 02
67 80 00 00 13 01 01 FE 23 2E 81 00 13 04 01 02
23 26 A4 FE 83 27 C4 FE 93 A7 57 00 13 F7 F7 0F
B7 17 40 00 93 87 07 80 23 A2 E7 00 13 00 00 00
03 24 C1 01 13 01 01 02 67 80 00 00 13 01 01 FE
23 2E 81 00 13 04 01 02 23 26 A4 FE B7 17 40 00
93 87 07 80 03 27 C4 FE 13 77 67 00 23 A4 E7 00
13 00 00 00 03 24 C1 01 13 01 01 02 67 80 00 00
13 01 01 FE 23 2E 81 00 13 04 01 02 23 26 A4 FE
83 27 C4 FE 93 E7 A7 01 23 26 F4 FE 03 27 C4 FE
93 07 E0 01 63 1A F7 00 B7 17 40 00 93 87 07 80
13 07 10 00 23 A6 E7 00 13 00 00 00 03 24 C1 01
13 01 01 02 67 80 00 00 13 01 01 FE 23 2E 81 00
13 04 01 02 23 26 A4 FE B7 17 40 00 93 87 07 80
03 27 C4 FE 13 47 A7 02 23 A8 E7 00 13 00 00 00
03 24 C1 01 13 01 01 02 67 80 00 00 13 01 01 FE
23 2E 81 00 13 04 01 02 23 26 A4 FE 83 27 C4 FE
93 97 37 00 23 26 F4 FE 03 27 C4 FE 93 07 00 04
63 1A F7 00 B7 17 40 00 93 87 07 80 13 07 10 00
23 AA E7 00 13 00 00 00 03 24 C1 01 13 01 01 02
67 80 00 00 13 01 01 FE 23 2E 81 00 13 04 01 02
23 26 A4 FE B7 17 04 00 93 87 07 E0 03 27 C4 FE
13 57 C7 00 23 AC E7 00 13 00 00 00 03 24 C1 01
13 01 01 02 67 80 00 00 13 01 01 FE 23 2E 81 00
13 04 01 02 23 26 A4 FE 83 27 C4 FE 93 D7 37 40
23 26 F4 FE 03 27 C4 FE 93 07 00 C0 63 1A F7 00
B7 17 40 00 93 87 07 80 13 07 10 00 23 AE E7 00
13 00 00 00 03 24 C1 01 13 01 01 02 67 80 00 00
13 01 01 FE 23 2E 81 00 13 04 01 02 23 26 A4 FE
23 24 B4 FE 03 27 C4 FE 83 27 84 FE B3 07 F7 00
23 26 F4 FE 03 27 C4 FE 93 07 30 24 63 1A F7 00
B7 17 40 00 93 87 07 80 13 07 10 00 23 A0 E7 02
13 00 00 00 03 24 C1 01 13 01 01 02 67 80 00 00
13 01 01 FE 23 2E 81 00 13 04 01 02 23 26 A4 FE
23 24 B4 FE 03 27 C4 FE 83 27 84 FE B3 27 F7 00
13 F7 F7 0F B7 17 40 00 93 87 07 80 23 A2 E7 02
13 00 00 00 03 24 C1 01 13 01 01 02 67 80 00 00
13 01 01 FE 23 2E 81 00 13 04 01 02 23 26 A4 FE
83 27 C4 FE B3 37 F0 00 13 F7 F7 0F B7 17 40 00
93 87 07 80 23 A4 E7 02 13 00 00 00 03 24 C1 01
13 01 01 02 67 80 00 00 13 01 01 FE 23 2E 81 00
13 04 01 02 23 26 A4 FE 23 24 B4 FE B7 17 40 00
93 87 07 80 83 26 C4 FE 03 27 84 FE 33 F7 E6 00
23 A6 E7 02 13 00 00 00 03 24 C1 01 13 01 01 02
67 80 00 00 13 01 01 FE 23 2E 81 00 13 04 01 02
23 26 A4 FE 23 24 B4 FE 03 27 C4 FE 83 27 84 FE
B3 67 F7 00 23 26 F4 FE 03 27 C4 FE B7 17 00 00
93 87 67 ED 63 1A F7 00 B7 17 40 00 93 87 07 80
13 07 10 00 23 A8 E7 02 13 00 00 00 03 24 C1 01
13 01 01 02 67 80 00 00 13 01 01 FE 23 2E 81 00
13 04 01 02 23 26 A4 FE 23 24 B4 FE B7 17 40 00
93 87 07 80 83 26 C4 FE 03 27 84 FE 33 C7 E6 00
23 AA E7 02 13 00 00 00 03 24 C1 01 13 01 01 02
67 80 00 00 13 01 01 FE 23 2E 81 00 13 04 01 02
23 26 A4 FE 23 24 B4 FE 83 27 84 FE 03 27 C4 FE
B3 17 F7 00 23 26 F4 FE 03 27 C4 FE B7 87 00 00
63 1A F7 00 B7 17 40 00 93 87 07 80 13 07 10 00
23 AC E7 02 13 00 00 00 03 24 C1 01 13 01 01 02
67 80 00 00 13 01 01 FE 23 2E 81 00 13 04 01 02
23 26 A4 FE 23 24 B4 FE B7 17 04 00 93 87 07 E0
03 27 84 FE 83 26 C4 FE 33 D7 E6 00 23 AE E7 02
13 00 00 00 03 24 C1 01 13 01 01 02 67 80 00 00
13 01 01 FE 23 2E 81 00 13 04 01 02 23 26 A4 FE
23 24 B4 FE B7 17 40 00 93 87 07 80 83 26 84 FE
03 27 C4 FE 33 87 E6 40 23 A0 E7 04 13 00 00 00
03 24 C1 01 13 01 01 02 67 80 00 00 13 01 01 FE
23 2E 81 00 13 04 01 02 23 26 A4 FE 23 24 B4 FE
83 27 84 FE 03 27 C4 FE B3 57 F7 40 23 26 F4 FE
03 27 C4 FE 93 07 00 C0 63 1A F7 00 B7 17 40 00
93 87 07 80 13 07 10 00 23 A2 E7 04 13 00 00 00
03 24 C1 01 13 01 01 02 67 80 00 00 13 01 01 FE
23 2E 81 00 13 04 01 02 23 26 A4 FE 23 24 B4 FE
03 27 C4 FE 83 27 84 FE 63 0A F7 00 B7 17 40 00
93 87 07 80 13 07 10 00 23 A4 E7 04 13 00 00 00
03 24 C1 01 13 01 01 02 67 80 00 00 13 01 01 FE
23 2E 81 00 13 04 01 02 23 26 A4 FE 23 24 B4 FE
03 27 C4 FE 83 27 84 FE 63 1A F7 00 B7 17 40 00
93 87 07 80 13 07 10 00 23 A6 E7 04 13 00 00 00
03 24 C1 01 13 01 01 02 67 80 00 00 13 01 01 FE
23 2E 81 00 13 04 01 02 23 26 A4 FE 23 24 B4 FE
03 27 C4 FE 83 27 84 FE 63 4A F7 00 B7 17 40 00
93 87 07 80 13 07 10 00 23 A8 E7 04 13 00 00 00
03 24 C1 01 13 01 01 02 67 80 00 00 13 01 01 FE
23 2E 81 00 13 04 01 02 23 26 A4 FE 23 24 B4 FE
03 27 C4 FE 83 27 84 FE 63 5A F7 00 B7 17 40 00
93 87 07 80 13 07 10 00 23 AA E7 04 13 00 00 00
03 24 C1 01 13 01 01 02 67 80 00 00 13 01 01 FF
23 26 11 00 23 24 81 00 13 04 01 01 13 05 00 00
EF F0 1F A6 13 05 10 00 EF F0 DF A8 13 05 10 00
EF F0 DF AB 13 05 C0 00 EF F0 9F AE 13 05 90 02
EF F0 9F B2 13 05 80 00 EF F0 5F B5 37 15 00 00
EF F0 5F B9 37 F5 FF FF EF F0 1F BC 93 05 80 1C
13 05 B0 07 EF F0 DF BF 93 05 B0 0A 13 05 50 05
EF F0 9F CB B7 17 00 00 93 85 67 E4 13 05 20 4D
EF F0 5F CE 93 05 90 02 13 05 A0 02 EF F0 DF D2
93 05 30 00 37 15 00 00 EF F0 DF D5 93 05 C0 00
37 15 00 00 EF F0 1F DA 93 05 A0 07 13 05 B0 07
EF F0 1F DD 93 05 30 00 37 F5 FF FF EF F0 1F E0
93 05 90 00 13 05 50 00 EF F0 5F E4 93 05 A0 02
13 05 A0 02 EF F0 9F E7 93 05 40 00 13 05 90 00
EF F0 DF EA 93 05 70 00 13 05 10 00 EF F0 1F EE
13 00 00 00 13 85 07 00 83 20 C1 00 03 24 81 00
13 01 01 01 67 80 00 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 17 01 40 00 13 01 41 7B 13 05 00 00
93 05 00 00 EF F0 9F EB 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00
