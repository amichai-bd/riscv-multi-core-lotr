//place holder - see gpc_4t_log_gen.sv as reference
